module mario(ix,iy,oR,oG,oB,mask,clk);
input clk;
input [10:0] ix;
input [10:0] iy;
output [7:0] oR;
output [7:0] oG;
output [7:0] oB;
output mask;
reg [104:0] mario_r;
reg [104:0] mario_g;
reg [104:0] mario_b;
reg [26:0] mario_a;
parameter x_size = 26,y_size = 32;
wire mask;

assign oR = (ix<x_size&&iy<y_size)?{mario_r[4*ix+3],mario_r[4*ix+2],mario_r[4*ix+1],mario_r[4*ix],4'b0000}:{ix[7:0]};
assign oG = (ix<x_size&&iy<y_size)?{mario_g[4*ix+3],mario_g[4*ix+2],mario_g[4*ix+1],mario_g[4*ix],4'b0000}:{iy[7:0]};
assign oB = (ix<x_size&&iy<y_size)?{mario_b[4*ix+3],mario_b[4*ix+2],mario_b[4*ix+1],mario_b[4*ix],4'b0000}:{ix+iy}; 
assign mask = (ix<x_size&&iy<y_size)?{mario_a[ix]}:0; 
always @(posedge clk)
begin
case(iy[5:0])
6'd0:mario_r=104'h000000feeffffff00000000000;
6'd1:mario_r=104'h000008defffffff00000000000;
6'd2:mario_r=104'h0000fbdeffffffff0000000000;
6'd3:mario_r=104'h0000acdeffffffeeffed000000;
6'd4:mario_r=104'h0000bcdeffffffffec98000000;
6'd5:mario_r=104'h000abcdefffffedca888000000;
6'd6:mario_r=104'h000aacdefffeec988880000000;
6'd7:mario_r=104'h009aabddedccdebba8ff000000;
6'd8:mario_r=104'hfaaaaabbb9adffb9efffff0000;
6'd9:mario_r=104'haaa999abb779dfc8cfffff0000;
6'd10:mario_r=104'hbaa999cfea77cfb56adfff0000;
6'd11:mario_r=104'hbba999dfeebaefe5138cef0000;
6'd12:mario_r=104'hfbba86afeefffffe8223c00000;
6'd13:mario_r=104'h0aba767addeefeeeeb21000000;
6'd14:mario_r=104'h00dc987679bddddeee0cdeff00;
6'd15:mario_r=104'hcdeffedcba977acddedddeffff;
6'd16:mario_r=104'hacdefffffffe92467cccedbeff;
6'd17:mario_r=104'h99bbeefddddee93657abdc9cee;
6'd18:mario_r=104'h9999bbcbaaaceb4ad357ad99cd;
6'd19:mario_r=104'h9988aaba689b9414922679979a;
6'd20:mario_r=104'h09988aba01221111111477bca8;
6'd21:mario_r=104'h000a986200000111111118bb99;
6'd22:mario_r=104'h0000754200000011111117987b;
6'd23:mario_r=104'h0000754100000001111116868a;
6'd24:mario_r=104'h0000743100000000001116667b;
6'd25:mario_r=104'h00005430000000000000156670;
6'd26:mario_r=104'h00095530000000000000155690;
6'd27:mario_r=104'h00084530000000000000355800;
6'd28:mario_r=104'h00865651000000000002457f00;
6'd29:mario_r=104'h00955674000100000004558000;
6'd30:mario_r=104'h00956787500000000000050000;
6'd31:mario_r=104'h00a56788a00000000000000000;
endcase
case(iy[5:0])
6'd0:mario_g=104'h00000001111115f00000000000;
6'd1:mario_g=104'h00000011111225c00000000000;
6'd2:mario_g=104'h00000111111223880000000000;
6'd3:mario_g=104'h00002111112222691111000000;
6'd4:mario_g=104'h00001111112221111111000000;
6'd5:mario_g=104'h00011111111111111111000000;
6'd6:mario_g=104'h00011111111112431110000000;
6'd7:mario_g=104'h002111111123689842ff000000;
6'd8:mario_g=104'h011111111137bdb9caceff0000;
6'd9:mario_g=104'h1111113652239ec899bdee0000;
6'd10:mario_g=104'h1111128ca6228ea4468acc0000;
6'd11:mario_g=104'h1111129daa75bec30158ab0000;
6'd12:mario_g=104'h0111116ddccbccca5101900000;
6'd13:mario_g=104'h00111126aa899a9aa810000000;
6'd14:mario_g=104'h00eb6531235667789a0cdfff00;
6'd15:mario_g=104'hdefffed51123345687cdefffff;
6'd16:mario_g=104'hbdeffffe42212332229deedfff;
6'd17:mario_g=104'habcdfffe51111257649bedbeff;
6'd18:mario_g=104'haabbdcdb3111125be669ceabde;
6'd19:mario_g=104'hbaaabbc921112446a5579aa8ab;
6'd20:mario_g=104'h0ba99bcb322344444446976665;
6'd21:mario_g=104'h000ba841333344444455356645;
6'd22:mario_g=104'h00003211333344445555445446;
6'd23:mario_g=104'h00004221333333444555444346;
6'd24:mario_g=104'h00004222233333334444433347;
6'd25:mario_g=104'h00003222233333333344433350;
6'd26:mario_g=104'h00052233222223333333332360;
6'd27:mario_g=104'h00052233333333333333323500;
6'd28:mario_g=104'h00532333333332000433324000;
6'd29:mario_g=104'h00632343333300000053336000;
6'd30:mario_g=104'h00623444400000000000000000;
6'd31:mario_g=104'h00523445500000000000000000;
endcase
case(iy[5:0])
6'd0:mario_b=104'h00000001111115f00000000000;
6'd1:mario_b=104'h00000011111115c00000000000;
6'd2:mario_b=104'h00000111111113880000000000;
6'd3:mario_b=104'h00002111111122691111000000;
6'd4:mario_b=104'h00001111111111111111000000;
6'd5:mario_b=104'h00011111111111111111000000;
6'd6:mario_b=104'h00011111111112321110000000;
6'd7:mario_b=104'h002111111113468732ff000000;
6'd8:mario_b=104'h0111111111159ab9989bcc0000;
6'd9:mario_b=104'h1111112440017bb9778abb0000;
6'd10:mario_b=104'h1111126984006b833568990000;
6'd11:mario_b=104'h1111127a77538a920146780000;
6'd12:mario_b=104'h0111104aa99899974101600000;
6'd13:mario_b=104'h00110004776677777610000000;
6'd14:mario_b=104'h00fb642011345556780cefff00;
6'd15:mario_b=104'heffffed51013334466deefffff;
6'd16:mario_b=104'hceffffff41123884329dffefff;
6'd17:mario_b=104'hccdefffe511114ba978cfeceff;
6'd18:mario_b=104'hccccedec411114976b99debcde;
6'd19:mario_b=104'hccbcdcda41114ac85cb8aba8ac;
6'd20:mario_b=104'h0ccbbcdca779bcdcbccb963223;
6'd21:mario_b=104'h000db943a99abcccdddd922222;
6'd22:mario_b=104'h00002103999abbcddeeda22113;
6'd23:mario_b=104'h000021139999abccddddb21123;
6'd24:mario_b=104'h000021357a999aabbcccc21124;
6'd25:mario_b=104'h0000104778999999aabba21120;
6'd26:mario_b=104'h000311488888899aa9aa821140;
6'd27:mario_b=104'h000311489988889aaaa9511200;
6'd28:mario_b=104'h0022112799a99a000ba8312000;
6'd29:mario_b=104'h0031111499aaf00000a4113000;
6'd30:mario_b=104'h00311112400000000000000000;
6'd31:mario_b=104'h00511112000000000000000000;
endcase
case(iy[5:0])
6'd0:mario_a=26'b00000000011110000000000000;
6'd1:mario_a=26'b00000001111111000000000000;
6'd2:mario_a=26'b00000011111111100000000000;
6'd3:mario_a=26'b00000111111111100000000000;
6'd4:mario_a=26'b00000111111111111110000000;
6'd5:mario_a=26'b00001111111111111110000000;
6'd6:mario_a=26'b00001111111111111100000000;
6'd7:mario_a=26'b00011111111111110000000000;
6'd8:mario_a=26'b00011111111111110011100000;
6'd9:mario_a=26'b00111111111111111111100000;
6'd10:mario_a=26'b01111111111111111111100000;
6'd11:mario_a=26'b01111111111111111111100000;
6'd12:mario_a=26'b00111111111111111110000000;
6'd13:mario_a=26'b00011111111111111100000000;
6'd14:mario_a=26'b00001111111111111000000000;
6'd15:mario_a=26'b00111111111111111001111100;
6'd16:mario_a=26'b11111111111111111111111110;
6'd17:mario_a=26'b11111111111111111111111110;
6'd18:mario_a=26'b11111111111111111111111110;
6'd19:mario_a=26'b01111111111111111111111110;
6'd20:mario_a=26'b00011110111111111110011110;
6'd21:mario_a=26'b00001100111111111111011111;
6'd22:mario_a=26'b00000111111111111111111111;
6'd23:mario_a=26'b00000111111111111111111110;
6'd24:mario_a=26'b00000111111111111111111110;
6'd25:mario_a=26'b00001111111111111111111100;
6'd26:mario_a=26'b00001111111111111111111100;
6'd27:mario_a=26'b00001111111111001111111000;
6'd28:mario_a=26'b00011111111100000001111000;
6'd29:mario_a=26'b00011111100000000000110000;
6'd30:mario_a=26'b00011110000000000000000000;
6'd31:mario_a=26'b00001110000000000000000000;
endcase
end
endmodule
