module arrow(ix,iy,mask,clk);
input clk;
input [10:0] ix;
input [10:0] iy;
output mask;

reg [64:0] arrow_a;
parameter x_size = 64,y_size = 64;
wire mask;
assign mask = (ix<x_size&&iy<y_size)?{arrow_a[ix[5:0]]}:0; 
always @(posedge clk)
begin
case(iy[5:0])
7'd0:arrow_a=64'b0000000000000000000000000000000000000000000000000000000000000000;
7'd1:arrow_a=64'b0000000000000000000000000001111111111000000000000000000000000000;
7'd2:arrow_a=64'b0000000000000000000000111111111111111111110000000000000000000000;
7'd3:arrow_a=64'b0000000000000000000011111111111111111111111100000000000000000000;
7'd4:arrow_a=64'b0000000000000000001111111111111111111111111111000000000000000000;
7'd5:arrow_a=64'b0000000000000000111111111111111111111111111111110000000000000000;
7'd6:arrow_a=64'b0000000000000011111111111111111111111111111111111100000000000000;
7'd7:arrow_a=64'b0000000000000111111111111111111111111111111111111110000000000000;
7'd8:arrow_a=64'b0000000000001111111111111111111111111111111111111111000000000000;
7'd9 :arrow_a=64'b0000000000011111111111111111111111111111111111111111100000000000;
7'd10:arrow_a=64'b0000000000111111111111111111111111111111111111111111110000000000;
7'd11:arrow_a=64'b0000000001111111111111111111111111001111111111111111111000000000;
7'd12:arrow_a=64'b0000000011111111111111111111111110000011111111111111111100000000;
7'd13:arrow_a=64'b0000000111111111111111111111111100000001111111111111111110000000;
7'd14:arrow_a=64'b0000001111111111111111111111111100000000111111111111111111000000;
7'd15:arrow_a=64'b0000001111111111111111111111111100000000011111111111111111000000;
7'd16:arrow_a=64'b0000011111111111111111111111111110000000001111111111111111100000;
7'd17:arrow_a=64'b0000011111111111111111111111111111000000000111111111111111100000;
7'd18:arrow_a=64'b0000111111111111111111111111111111100000000011111111111111110000;
7'd19:arrow_a=64'b0000111111111111111111111111111111110000000001111111111111110000;
7'd20:arrow_a=64'b0001111111111111111111111111111111111000000000111111111111111000;
7'd21:arrow_a=64'b0001111111111111111111111111111111111100000000001111111111111000;
7'd22:arrow_a=64'b0011111111111111111111111111111111111110000000000111111111111100;
7'd23:arrow_a=64'b0011111111111111111111111111111111111111000000000011111111111100;
7'd24:arrow_a=64'b0011111111111111111111111111111111111111100000000001111111111100;
7'd25:arrow_a=64'b0011111111111111111111111111111111111111110000000000111111111100;
7'd26:arrow_a=64'b0011111111111111111111111111111111111111111000000000011111111100;
7'd27:arrow_a=64'b0111111111111111111111111111111111111111111110000000001111111110;
7'd28:arrow_a=64'b0111111111111111111111111111111111111111111110000000000111111110;
7'd29:arrow_a=64'b0111111111000000000000000000000000000000000000000000000011111110;
7'd30:arrow_a=64'b0111111110000000000000000000000000000000000000000000000001111110;
7'd31:arrow_a=64'b0111111110000000000000000000000000000000000000000000000001111110;
7'd32:arrow_a=64'b0111111110000000000000000000000000000000000000000000000001111110;
7'd33:arrow_a=64'b0111111110000000000000000000000000000000000000000000000001111110;
7'd34:arrow_a=64'b0111111111000000000000000000000000000000000000000000000011111110;
7'd35:arrow_a=64'b0111111111111111111111111111111111111111111110000000000111111110;
7'd36:arrow_a=64'b0111111111111111111111111111111111111111111100000000001111111110;
7'd37:arrow_a=64'b0011111111111111111111111111111111111111111000000000011111111100;
7'd38:arrow_a=64'b0011111111111111111111111111111111111111110000000000111111111100;
7'd39:arrow_a=64'b0011111111111111111111111111111111111111100000000001111111111100;
7'd40:arrow_a=64'b0011111111111111111111111111111111111111000000000011111111111100;
7'd41:arrow_a=64'b0011111111111111111111111111111111111110000000001111111111111000;
7'd42:arrow_a=64'b0001111111111111111111111111111111111100000000011111111111111000;
7'd43:arrow_a=64'b0001111111111111111111111111111111111000000000111111111111111000;
7'd44:arrow_a=64'b0000111111111111111111111111111111110000000001111111111111110000;
7'd45:arrow_a=64'b0000111111111111111111111111111111100000000011111111111111110000;
7'd46:arrow_a=64'b0000011111111111111111111111111111000000000111111111111111100000;
7'd47:arrow_a=64'b0000011111111111111111111111111110000000001111111111111111100000;
7'd48:arrow_a=64'b0000001111111111111111111111111100000000011111111111111111000000;
7'd49:arrow_a=64'b0000001111111111111111111111111100000000111111111111111111000000;
7'd50:arrow_a=64'b0000000111111111111111111111111100000001111111111111111110000000;
7'd51:arrow_a=64'b0000000011111111111111111111111110000011111111111111111100000000;
7'd52:arrow_a=64'b0000000001111111111111111111111111111111111111111111111000000000;
7'd53:arrow_a=64'b0000000000111111111111111111111111111111111111111111110000000000;
7'd54:arrow_a=64'b0000000000011111111111111111111111111111111111111111100000000000;
7'd55:arrow_a=64'b0000000000001111111111111111111111111111111111111111000000000000;
7'd56:arrow_a=64'b0000000000000111111111111111111111111111111111111110000000000000;
7'd57:arrow_a=64'b0000000000000011111111111111111111111111111111111100000000000000;
7'd58:arrow_a=64'b0000000000000000111111111111111111111111111111110000000000000000;
7'd59:arrow_a=64'b0000000000000000001111111111111111111111111111000000000000000000;
7'd60:arrow_a=64'b0000000000000000000011111111111111111111111100000000000000000000;
7'd61:arrow_a=64'b0000000000000000000000111111111111111111100000000000000000000000;
7'd62:arrow_a=64'b0000000000000000000000000001111111111000000000000000000000000000;
7'd63:arrow_a=64'b0000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule
