// --------------------------------------------------------------------
// Copyright (c) 2007 by Terasic Technologies Inc. 
// --------------------------------------------------------------------
//
// Permission:
//
//   Terasic grants permission to use and modify this code for use
//   in synthesis for all Terasic Development Boards and Altera Development 
//   Kits made by Terasic.  Other use of this code, including the selling 
//   ,duplication, or modification of any portion is strictly prohibited.
//
// Disclaimer:
//
//   This VHDL/Verilog or C/C++ source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  Terasic provides no warranty regarding the use 
//   or functionality of this code.
//
// --------------------------------------------------------------------
//           
//                     Terasic Technologies Inc
//                     356 Fu-Shin E. Rd Sec. 1. JhuBei City,
//                     HsinChu County, Taiwan
//                     302
//
//                     web: http://www.terasic.com/
//                     email: support@terasic.com
//
// --------------------------------------------------------------------
//
// Major Functions:	DE2 LTM module Timing control and output image data
//					form sdram 
//
// --------------------------------------------------------------------
//
// Revision History :
// --------------------------------------------------------------------
//   Ver  :| Author            		:| Mod. Date :| Changes Made:
//   V1.0 :| Johnny Fan				:| 07/06/30  :| Initial Revision
// --------------------------------------------------------------------

module ltp_controller(
						iCLK, 				// LCD display clock
						iRST_n, 			// systen reset
						// SDRAM SIDE 
						iREAD_DATA1, 		// R and G  color data form sdram 	
						iREAD_DATA2,		// B color data form sdram
						oREAD_SDRAM_EN,		// read sdram data control signal
						//LCD SIDE
						oHD,				// LCD Horizontal sync 
						oVD,				// LCD Vertical sync 	
						oDEN,				// LCD Data Enable
						oLCD_R,				// LCD Red color data 
						oLCD_G,             // LCD Green color data  
						oLCD_B,             // LCD Blue color data  
						);
//============================================================================
// PARAMETER declarations
//============================================================================
parameter H_LINE = 1056; 
parameter V_LINE = 525;
parameter Hsync_Blank = 46;   //H_SYNC + H_Back_Porch
parameter Hsync_Front_Porch = 210;
parameter Vertical_Back_Porch = 23; //V_SYNC + V_BACK_PORCH
parameter Vertical_Front_Porch = 22;
//===========================================================================
// PORT declarations
//===========================================================================
input			iCLK;   
input			iRST_n;
input	[15:0]	iREAD_DATA1;
input	[15:0]	iREAD_DATA2;
output			oREAD_SDRAM_EN;
output	[7:0]	oLCD_R;		
output  [7:0]	oLCD_G;
output  [7:0]	oLCD_B;
output			oHD;
output			oVD;
output			oDEN;
//=============================================================================
// REG/WIRE declarations
//=============================================================================
reg		[10:0]  x_cnt;  
reg		[9:0]	y_cnt; 
wire	[7:0]	read_red;
wire	[7:0]	read_green;
wire	[7:0]	read_blue; 
wire			display_area;
wire			oREAD_SDRAM_EN;
reg				mhd;
reg				mvd;
reg				mden;
reg				oHD;
reg				oVD;
reg				oDEN;
reg		[7:0]	oLCD_R;
reg		[7:0]	oLCD_G;	
reg		[7:0]	oLCD_B;
		
reg [7:0] time_count;
reg [15:0] distance;




reg	[7:0]	frame_count;

reg [9:0] move_x;
reg [9:0] move_y;

reg [956:0] marior,mariog,mariob;
wire [3:0] pixelr,pixelg,pixelb;
assign pixelr = {marior[4*(x_cnt-move_x)],marior[4*(x_cnt-move_x)+1],marior[4*(x_cnt-move_x)+2],marior[4*(x_cnt-move_x)+3]};
assign pixelg = {mariog[4*(x_cnt-move_x)],mariog[4*(x_cnt-move_x)+1],mariog[4*(x_cnt-move_x)+2],mariog[4*(x_cnt-move_x)+3]};
assign pixelb = {mariob[4*(x_cnt-move_x)],mariob[4*(x_cnt-move_x)+1],mariob[4*(x_cnt-move_x)+2],mariob[4*(x_cnt-move_x)+3]};
//assign pixel = marior[(x_cnt-move_x)];

parameter move_size_x = 239;
parameter move_size_y = 500;
assign	road1	  =  ((x_cnt>40 && x_cnt<150)  ) ? 1'b1: 1'b0;
assign	road2   =  ((x_cnt>750 && x_cnt<850 ) ) ? 1'b1: 1'b0;


//=============================================================================
// Structural coding
//=============================================================================

// This signal control reading data form SDRAM , if high read color data form sdram  .
assign	oREAD_SDRAM_EN = (	(x_cnt>Hsync_Blank-2)&& //214
							(x_cnt<(H_LINE-Hsync_Front_Porch-1))&& //1015
							(y_cnt>(Vertical_Back_Porch-1))&& // //34
							(y_cnt<(V_LINE - Vertical_Front_Porch)) //515
						 )?  1'b1 : 1'b0;
						
// This signal indicate the lcd display area .
assign	display_area = ((x_cnt>(Hsync_Blank-1)&& //>215
						(x_cnt<(H_LINE-Hsync_Front_Porch))&& //< 1016
						(y_cnt>(Vertical_Back_Porch-1))&& 
						(y_cnt<(V_LINE - Vertical_Front_Porch-1))
						))  ? 1'b1 : 1'b0;

assign	read_red 	= display_area ? iREAD_DATA2[9:2] : 8'b0;
assign	read_green 	= display_area ? {iREAD_DATA1[14:10],iREAD_DATA2[14:12]}: 8'b0;
assign	read_blue 	= display_area ? iREAD_DATA1[9:2] : 8'b0;

assign draw_circle = (x_cnt-300)*(x_cnt-300)+(y_cnt-300)*(y_cnt-300) < 40000 ? 1'b1:1'b0;


///////////////////////// x  y counter  and lcd hd generator //////////////////
always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
		begin
			x_cnt <= 11'd0;	
			mhd  <= 1'd0;  	
		end	
		else if (x_cnt == (H_LINE-1))
		begin
			x_cnt <= 11'd0;
			mhd  <= 1'd0;
		end	   
		else
		begin
			x_cnt <= x_cnt + 11'd1;
			mhd  <= 1'd1;
		end	
	end

always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
		begin
			y_cnt <= 10'd0;
			
			
			//frame_count <= 8'b0;
			move_x <= 0;
			move_y <= 0;
		end
		else if (x_cnt == (H_LINE-1))
		begin
			if (y_cnt == (V_LINE-1))
			begin
				y_cnt <= 10'd0;
				time_count <= time_count + 1;
			end
			else
			begin
				y_cnt <= y_cnt + 10'd1;	
				//frame_count <= (frame_count > 60)?  0 : frame_count+1;
			end
			
				
		end else if(x_cnt == 0&&y_cnt == (V_LINE-1))
		begin
			//move_x <= move_x+1;
			//move_y <= move_y+2;
		end
	end
////////////////////////////// touch panel timing //////////////////

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			mvd  <= 1'b1;
		else if (y_cnt == 10'd0)
			mvd  <= 1'b0;
		else
			mvd  <= 1'b1;
	end			

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			mden  <= 1'b0;
		else if (display_area)
			mden  <= 1'b1;
		else
			mden  <= 1'b0;
	end			

always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
			begin
				oHD	<= 1'd0;
				oVD	<= 1'd0;
				oDEN <= 1'd0;
				oLCD_R <= 8'd0;
				oLCD_G <= 8'd0;
				oLCD_B <= 8'd0;
			end
			

		else if 	((move_x<x_cnt && (x_cnt<move_x+move_size_x) && move_y<y_cnt && (y_cnt<move_y+move_size_y)) )
		begin
                oLCD_R	<= {pixelr,4'b0000};
                oLCD_G	<= {pixelg,4'b0000};
					 oLCD_B	<= {pixelb,4'b0000};
		end

		else
			begin
				oHD	<= mhd;
				oVD	<= mvd;
				oDEN <= mden;
				distance <= (x_cnt-300)*(x_cnt-300)+(y_cnt-300)*(y_cnt-300);
				oLCD_R <= draw_circle?time_count+(x_cnt-300)+(y_cnt-300):read_red;
				oLCD_G <= draw_circle?time_count+x_cnt:read_green;
				oLCD_B <= draw_circle?time_count+distance[15:8]:read_blue;
				//oLCD_R	<= {pixel,4'b0000};
            //oLCD_G	<= {8'hff};
				//oLCD_B	<= {8'hff};
			end		
	end
						
						
always@(posedge iCLK or negedge iRST_n)
begin
	case((y_cnt-move_y))
 
 10'd0:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd1:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd2:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeffeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd3:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeefeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd4:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd5:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd6:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd7:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd8:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd9:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd10:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd11:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd12:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffefefffeeefefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd13:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedccccccccdeffffeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd14:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeccdeffffffdedcceffffeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd15:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffecdfffffffffedefffdcdfffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd16:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffddffffffffffddedeffffddeffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd17:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffddeffffffffffedeeedfffffeceffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd18:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffddffffffffffffdeddedeffffffceffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd19:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffdedeffffffffffeeedddedfffffffddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd20:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffdffdddffffffffedfddddeedfffffffdefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd21:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffdffeeeeefffffffdeedddddeddfffffffdfeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd22:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffdefededefefffffeeeeddddddedfffffffeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd23:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffeeffededdffefffedededddddddedffffffedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd24:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffedfffededdeefeefddededddddddeddffffffeeeddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeeedeedeeedddddefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd25:marior=956'hffffffffffffffffffffffffffffffffffffffffffffefdffffeedddeeeeededddddccdddddedfffffffeeedeeeeeeeeeeeeeeeeeeeedeeeeeeeeeedeeeddeeddeddeddeeddddeddddddeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd26:marior=956'hfffffffffffffffffffffffffffffffffffffffffffefeefffeeedededddeeedddddbccdddddedffffffeeedeeeeeeeeeeeeeeeeeeeeedeededeedededddddededdddddddddedddddddddefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd27:marior=956'hfffffffffffffffffffffffffffffffffffffffffeeefeffffdedddddddddedddddcddcdcdddddefffffeeeddeeeeeeeeeeedddeededdededeeddddddddddddddddddddddddddddddddddddffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd28:marior=956'hffffffffffffffffffffffffffffffffffffffeeeeefeefffededdddddddddddddccfecdddddcddefffffeeddddddedddededededddeddddddddddddddddddddddddddddddddddddddddddddfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd29:marior=956'hfffffffffffffffffffffffffffffffffffffffefeeedffffeddddcbcdddddddcdceffdccddccdddfffffeeddeddedededddddddeeededdddddddddddddddddddddddddddddddddddddddddddffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd30:marior=956'hffffffffffffffffffffffffffffffffffffeeeeeeefeffffeedddcccdddddddcdcfffecdddcdccedffffeeccdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd31:marior=956'hffffffffffffffffffffffffffffffffffffeeeeeeeeeffffdedddcefccdcdddccdffffccddcdccecefffeedcddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd32:marior=956'hfffffffffffffffffffffffffffffffffffeeeeeeeeeffffededddceffbccdcdccfffffdcdccccdcddfffeedcdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd33:marior=956'hfffffffffffffffffffffffffffffffffffeeeeeeeeeffffeddddcdfffeccdcdbdffffffcccdccccdedfffecbddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd34:marior=956'hffffffffffffffffffffffffffffffffffeeeeeeeeeeffffdddddccffffebcccbeffffffecccccccddcdffecbdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd35:marior=956'hffffffffffffffffffffffffffffffffffeeeeeeeefeffffddddddcfffffebbbcffffffffccccccdccccdeebbddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd36:marior=956'hfffffffffffffffffffffffffffffffffeeeeeeeeeeefffeddcddccfffffffbbeffffffffecbcccdccdccfebbdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd37:marior=956'hfffffffffffffffffffffffffffffffffeeeeeeeeeeefffdcddcdcdfffffffecffffffffffcbccdcbccacfdacddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd38:marior=956'hfffffffffffffffffffffffffffffffffeeeeeeeeeeefffddcddccdfffffffffffffffffffebbccbccaceec9cdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd39:marior=956'hffffffffffffffffffffffffffffffffeeeeeeeeeeeefffdddcddcdffffffffffffffffffffcbccbcbbefeb9dddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddceffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd40:marior=956'hffffffffffffffffffffffffffffffffeeeeeeeeeeeefffccddcdcdfffffffffffffffffeffeccbcbadefdaaddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd41:marior=956'hfffffffffffffffffffffffffffffffeeeeeeeeeedddffeddddcccdfffffffffffffffffffeecbbcacdfec9bdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd42:marior=956'hfffffffffffffffffffffffffffffffeeeeeeeeeedeeefedddcccbdffffffffffffffeeeeeeeebbacddfdaacdddddddddcddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd43:marior=956'hfffffffffffffffffffffffffffffffeeeeeeeeeeddeefdcdddccbdfffffffffffffeffeeeeeecbaddfec9bdccccdccddddddcdcddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd44:marior=956'hfffffffffffffffffffffffffffffffeeeeeeeeddddeeedcccddcbdffffffeeeeeeefeeeeeededbccefca9cddddddddcddccdddddddcdcdddddcdddddddddddddddddddddddddddddddddddddddccddddddddcdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd45:marior=956'hffffffffffffffffffffffffffffffeeeeeeeeedddddeedcdccccbdfffffefeeeeeeeeeeeeddeeddeedb9bddcccccccccccccccccccdddddccddddddddddddddddddddddddddddddddddcdddcccccccccccdddcefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd46:marior=956'hffffffffffffffffffffffffffffffeeeeeeeedddddddedabcccccdfeeeffeeeeeeeeddddeeeeeeeedb99ccccccccccccccccccccccccccccdcccdcdcddddddcdddddddddddddddcddcdccccccccccccccccdddcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd47:marior=956'hffffffffffffffffffffffffffffffeeeeeeeddddddddefdbabccadeeeeeeeeedddeeefeeeddddcddcaacddeeeedddccccccccccccccccccccccccccccccdcdccccccdcddcdddcddccccccccccccccccccccccdccffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd48:marior=956'hffffffffffffffffffffffffffffffeeeeedddddddddddeeecaabbdeeeeeeddddeeeeddccccddeeeefffffffffffffffffeeddcccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccdcdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd49:marior=956'hffffffffffffffffffffffffffffffeeeeeddddddddddccffedcaaceeeeddeffedcccddeffffffffffffffffffffffffffffffffedccbbccccccccccccccccccccccccccccccccccccccccccccccccccccccccccdceffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd50:marior=956'hffffffffffffffffffffffffffffffeeeeddddddddddddbcefeedbcddddeeedccdeeffffffffffffffffffffffffffffffffffffeffeedcbbbbcccccccccccccccccccccccccccccccccccccccccccccccccccccccbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd51:marior=956'hffffffffffffffffffffffffffffffeeeedddddddddddddbcefedddddeedccdefffffffffffffffffffffffffffffffffffffffffeeeeeeecbbbbbbccccccccccccccccccccccccccccccccccccccccccccccccccccdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd52:marior=956'hfffffffffffffffffffffffffffffeeeeddddddddddddddcabdffdcdedddeffffffffffffffffffffffffffffffffffffffffffffefeeeeeeedbbbbbbbbbbbcccccccccccccccccccccccccccccccccccccccccccccceffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd53:marior=956'hfffffffffffffffffffffffffffffeeeeddddddddddddddddbacdeeedefffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeedcbabbbbbbbbbbbcbccccccccccccccccccccccccccccccccccccccdeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd54:marior=956'hfffffffffffffffffffffffffffffeeeddddddddddddddddddbaaceffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeedcaaaabbbbbbbbbbbcbcccccccccccccccccccccccccccccccccccdeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd55:marior=956'hfffffffffffffffffffffffffffffeedddddddddddddddddcccdefffffffffffffffffffffeffeeeeeeeefefffffffffffffffffeeefefeeeeeeeeeeecaaaaabbbbbbbbbbbbbcbcccccccccccccccccccccccccccccccdeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd56:marior=956'hfffffffffffffffffffffffffffffeedddddddddddddddccdeffffffffffffffeeeeeddddddccdccdccdccccccdddddeeeeefffffefeeeeeeeeeeeeeeedbaaaaaaaabbbbbbbbbbbbbbcbcbcbbcbcbbbbbbbccccccccccddeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd57:marior=956'hfffffffffffffffffffffffffffffeddddddddddddddcdeffffffffffeeeedddddccccbbbbbaabaabaabaababbbbbbbccccdddeeeefffeeeeeeeeeeeeeeedb9aaaaaabbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbccccccccddddeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd58:marior=956'hfffffffffffffffffffffffffffffeeddddddddddccdeffffffffeeddddccbbbbbaa999999a999999999999999999aaaaaabbbbbccddeeeeeeeeeeeeeeeeeeda999aaaaaababbbbbbbbbbbbbbbbbbbbbbbbbbbbcbcccccddddddeefffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd59:marior=956'hfffffffffffffffffffffffffffffedddddddddddeffffffeeedddcccbba99999999999999999999999999999999999999999aaaabbbbccdeeeeeeeeeeeeeeeeca999999aaaaabbbbbbbbbbbbbbbbbbbbbbbbbbbbccccccdddddddeffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd60:marior=956'hfffffffffffffffffffffffffffffeddddddddeffffffeedcccbaaaa9a9999999999999999999999999999999999898989999999999aaaaabbcdeeeeeeeeeeeeedb9999999aaaaaabbbbbbbbbbbbbbbbbbbbbbbbbbbccccdddddddddfffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd61:marior=956'hfffffffffffffffffffffffffffffeddddddfffffeeddcbbaa999999999999999999999999999999999999999999898888888888999999aaaaaabccdeeeeeeeeeeeda99999999aaaaaaaaaabbbabbbbbbbbbbbbbbbbbccccdddddddddffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd62:marior=956'hfffffffffffffffffffffffffffffedddeffffedddcbaa99999999999999999999999999999999999999999999988888888888888888899999aaaaaabcddeeeedeeedb99999999aaaaaaaaaaabaaabbbbbbbbbbbbbbbbccccddddddddcfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd63:marior=956'hfffffffffffffffffffffffffffffddefffedcdccaa999999999999999999999999999999999999999999999988888888888888888888888899999aaaaabcdeeedddddca9999999aaaaaaaaaaaaaaaabbabbbbbbbbbbbccccccddddddcdffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd64:marior=956'hfffffffffffffffffffffffffffffefffddcbbaa9a9999999999999999999999999999999999999999998888888888888899999999988888888889999aaaaabcddedddddb99999999aaaaaaaaaaaaaaaaaaaabbbbbbbbbcccccccccdcdcdfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd65:marior=956'hffffffffffffffffffffffffffffffedccba9999999999999999999999999999999999999999998888888888888877766421122334456678888888889999aaaabbcddddddc999999999aaaaaaaaaaaaaaaaaaaabbbbbbbbccccccccccccbeffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd66:marior=956'hffffffffffffffffffffffffffffeddcbaa9999999999999999999999999999999999999888888878888888888888776300000000000000014677888889999aaaaabcdddddc9899999aaaaaaaaaaaaaaaaaaaaaaabbbbbbbbccccccccccccffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd67:marior=956'hffffffffffffffffffffffffffedcbba999999999999999999999999999999999999888777778888888888888888876100000000000000000036667778888899a9aaabbcdddca8999999aaaaaaaaaaaaaaaaaaaaaaabbbbbbbcbccccccccbdfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd68:marior=956'hfffffffffffffffffffffffffdccb999999999999999999999999999999999888887777888888888989999999988861000000011001000000004777777777888999aaaaabcddc98999999aaaaaaaaaaaaaaaaaaaaaaaabbbbbbbbbcccccccbfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd69:marior=956'hfffffffffffffffffffffffedcbaa999999999999999999999999999999988887777888888899999999999999998620001111111110101000001677888777777889999aaaabcdc9899999aaaaaaaaaaaaaaaaaaaaaaaaaabbbbbbbbbbbcccbcffffffffffffffffffffffffffffffffffffffffffffffff;
10'd70:marior=956'hffffffffffffffffffffffedba9999999999999999999999999998888888877788888899999999999999999999972011111111111111111100002788888888777778899aaaaabcca8999aaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbbbbbbbbbbbbefffffffffffffffffffffffffffffffffffffffffffffff;
10'd71:marior=956'hfffffffffffffffffffffdcaa999999999999999999999999988888888777788888999999999999999aaaaaa99830011111111111111111111000588888888888776788999aaaabba999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbbbbbbbbbbdfffffffffffffffffffffffffffffffffffffffffffffff;
10'd72:marior=956'hfffffffffffffffffffecba9999999999999999999999999988888887778888899999999999a9aaaaaaaaaaa996001111111111111111111111102888999888888877678899aaaaaa999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbabbbbfffffffffffffffffffffffffffffffffffffffffffffff;
10'd73:marior=956'hffffffffffffffffffecba9999999999999999999999998888888766788889999999999aaaaaaaaaaaaaaaaa982011111111111111111111111100699999999988888776788899aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbeffffffffffffffffffffffffffffffffffffffffffffff;
10'd74:marior=956'hfffffffffffffffffecba9999999999999999999999988888887666788899999999aaaaaaaaaaaaaaaaaaaaa95111111111111100000000111111039999999999998888877788899aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbadffffffffffffffffffffffffffffffffffffffffffffff;
10'd75:marior=956'hfffffffffffffffffcba9999999999999999999999888888886556778899999aaaaaaaaaaaaaaaaaaaaaaaaa920111111111001245555431001111189aaaaa9999999998887678889aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbacffffffffffffffffffffffffffffffffffffffffffffff;
10'd76:marior=956'hffffffffffffffffdb99999999999999999999998888888764100014789999aaaaaaaaaaaaaaaaababbbbbaa711111111002579aaaaaaaaa85201106aaaaaaaaaaaaaaa99998767888999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbbbffffffffffffffffffffffffffffffffffffffffffffff;
10'd77:marior=956'hfffffffffffffffeba9999999999999999999988888888762000000015899aaaaaaaaaaaaaaabbbbbbbbbbba401111110369aaaabbbbbbbbbba62004aaaaaaaaaaaaaaaaaaaa984467888999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbbefffffffffffffffffffffffffffffffffffffffffffff;
10'd78:marior=956'hfffffffffffffffca99999999999999999999988888877520111111000599aaaaaaaaaabbbbbbbbbbbbbbbb9211111016aabbbbbbbbbbbbbbbbba503aabbbbbbaabababbbbbbaa72334688899aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbadfffffffffffffffffffffffffffffffffffffffffffff;
10'd79:marior=956'hffffffffffffffeba99999999999999999999888888765201111111000059aaaaaaabbabbbbbbbbbbbbbbbb81111104abbbbbbbbbbbbbbbbbbbbbb729bbbbbbbbbbbbbbbbbbbbb9434334568899aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbacfffffffffffffffffffffffffffffffffffffffffffff;
10'd80:marior=956'hffffffffffffffca999999999999999999998888887753111111111111006aaaaabbbbbbbbbbbbbbbbbbbbb7011115bbbbbbbbbbbbbbbbbbbbbbbbb9abbbbbbbbbbbbbbbbbccbba63444444568999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbacfffffffffffffffffffffffffffffffffffffffffffff;
10'd81:marior=956'hffffffffffffffc99999999999999999999888888776421111111111111028aaaabbbbbbbbbbbbbbbbbbbbb501107bccccccccccccccbcccbbbbbbbccbbbbbbbbbbbbcccccccccb834444455456899aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbacfffffffffffffffffffffffffffffffffffffffffffff;
10'd82:marior=956'hfffffffffffffeb99999999999999999888888887765421111111111111104aabbbbbbbbbbbbbbbbbbbbbbb40117ccccccccccccccccccccccccccccccccccccccccccccccccccc94444555555556899aaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbacfffffffffffffffffffffffffffffffffffffffffffff;
10'd83:marior=956'hfffffffffffffea999999999999999998888888877654111111211111111119bbbbbbbbbbbbbbbbbccccccb4015bccccccccccccccccccccccccccccccccccccccccccccccccccca4445555555555579aaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbacfffffffffffffffffffffffffffffffffffffffffffff;
10'd84:marior=956'hfffffffffffffea999999999999999988888888776554111112222212111106abbbbbbbbbbbbccccccccccb404accccccccccccccccccccccccccccccccccccccccccccccccccccb54455555555555579aaaaaaaaaaaaaaaaaaaaaaaaaaaaabbacfffffffffffffffffffffffffffffffffffffffffffff;
10'd85:marior=956'hfffffffffffffea999999999999988888888888776573112222222222211102abbbbbbbbbcccccccccccccc419cccccccccccccccccccccccccccccccccccccccccccccccccccccb5445555555555555699999aaa9aa9999999999aaaaaaaabbacfffffffffffffffffffffffffffffffffffffffffffff;
10'd86:marior=956'hfffffffffffffea9999999999998988888888877765721122222222222211118bbbbbbccccccccccccccccc45ccccccccccbaabbbcccccccccccccccccddddddcdddccdccccccccc644555555555555556899999999998888998899aaaaaaabbacfffffffffffffffffffffffffffffffffffffffffffff;
10'd87:marior=956'hffffffffffffffb9999999999998888888888887766811221367888875321105bbbbccccccccccccccddddd7bddddddcbaaabbbbbbbbccddddddddddddddddddddddddddddddcccc645555555555555555689999989bdefffffedb989aaaaabbacfffffffffffffffffffffffffffffffffffffffffffff;
10'd88:marior=956'hffffffffffffffd99999999999988888888888777678111269aaaaaaaa974202accccccccccccddddeeeeeeeeeedddcaabcccccccccbbcdeeeefffffffffeeeeeeeedddddddddccc6455555555555555555689989dfffffffffffffda9aaaabbadfffffffffffffffffffffffffffffffffffffffffffff;
10'd89:marior=956'hfffffffffffffffa99999999999888888888887766871117aaaabbbbbbba95118ccccccccdddeeeefffffffffeeedcabcccdddddddddcbceffffffffffffffffffffffeeeeddddcc74555555555555556554677afffffffffffffffffc9aabbbbdfffffffffffffffffffffffffffffffffffffffffffff;
10'd90:marior=956'hfffffffffffffffd9999998989888888888888777698115aaabbbbbbbbbbba515cccccdddeeeffffffffffffffeecabcddddddddddddddccffffffffffffffffffffffffffeedddc7555555555555555655433bfffffffffffffffffffdaabbbbefffffffffffffffffffffffffffffffffffffffffffff;
10'd91:marior=956'hffffffffffffffffc99999988888888888888877769813aabbbbbbbbbcccccb63ccdddeeffffffffffffffffffedbbdddeeeeeeeeeeeeedcdffffffffffffffffffffffffffeeedd855555555555566566531bfffffffffffffffffffffeaabbbffffffffffffffffffffffffffffffffffffffffffffff;
10'd92:marior=956'hfffffffffffffffffb999998888888888888887776a917bbbbbbbbbccccccccb8bdeeeffffffffffffffffffffecbdeeeeeeeeeeffeeefedceffffffffffffffffffffffffffeedd856555555666565566527fffffffffffffffffffffffeabacffffffffffffffffffffffffffffffffffffffffffffff;
10'd93:marior=956'hffffffffffffffffffa99999898888888888887776a94abbbbbbbccccccccccccdeefffffffffffffffffffffedbceeeeeeeeffc7321249eddeffffffffffffffffffffffffffeed86665555556666666545effffffffffffffffffffffffcaadffffffffffffffffffffffffffffffffffffffffffffff;
10'd94:marior=956'hfffffffffffffffffffb9999998888888888887776aaabbbbbbbccccbbbbcccdeefffffffffffffffffffffffecbdeeeeeeefc4112222112bddffffffffffffffffffffffffffeed7666665566666666653affffffffffffffffffffffffffbaeffffffffffffffffffffffffffffffffffffffffffffff;
10'd95:marior=956'hffffffffffffffffffffc999989888888888888776abbbbbbbbccbbbaaababcdeffffffffffffffffffffffffecceeeeeeef9112222222211adeffffffffffffffffffffffffffec7666665566666666655dfffffffffffeeeeeefffffffffdbfffffffffffffffffffffffffffffffffffffffffffffff;
10'd96:marior=956'hfffffffffffffffffffffca9998888888888888877abbbbbbccccba9acccccbceffffffffffffffffffffffffdbdeeeeeefa12222222222212beffffffffffffffffffffffffffeb7776666666666666658efffffffffeeeeddddeeffffffffceffffffffffffffffffffffffffffffffffffffffffffff;
10'd97:marior=956'hffffffffffffffffffffffebaa9998988888888887acbbbbbcccbb9bcccccddccefffffffffffffffffffffffdbdeeeeefc2222222222222213dffffffffffffffffffffffffffea776666666666665665bffffffffeeeedddddddeefffffffdcffffffffffffffffffffffffffffffffffffffffffffff;
10'd98:marior=956'hffffffffffffffffffffffffdbaaaaa99999aaa987bcccccccccb9acccdddddeddfffffffffffffffffffffffccdeeeeef512222322222222207ffffffffffffffffffffffffffd8777666666666656666cfffffffeeedddddeeeeeefffffffebefffffffffffffffffffffffffffffffffffffffffffff;
10'd99:marior=956'hffffffffffffffffffffffffffecbabbbbbbbbbba8bdcccccccca8ccdddddefc97cffffffffffffffffffffffccdeeeeec222222323322222212cfffffffffffffffffffffffffb8877766666666666666dffffffeeddddeffffffffffffffffbcfffffffffffffffffffffffffffffffffffffffffffff;
10'd100:marior=956'hfffffffffffffffffffffffffffffeccbbbbbbbbcabdcccccccb9addddeeec31114effffffffffffffffffffecddeeeef71223333333222222219ffffffffffffffffffffffffe98887777666666666668dffffffedddeffffffffffffffffffdbeffffffffffffffffffffffffffffffffffffffffffff;
10'd101:marior=956'hffffffffffffffffffffffffffffffffffffffffffddcccccccb9cddeeefa2122219ffffffffffffffffffffecdddeeee41122233322222222217ffffffffffffffffffffffffd88888776666666566668dfffffedddffffffffffffffffffffebdffffffffffffffffffffffffffffffffffffffffffff;
10'd102:marior=956'hfffffffffffffffffffffffffffffffffffffffffffecccccccb9ddeeefb22222213ffffffffffffffffffffecdddeeed1111222228db32322215efffffffffffffffffffffffc88888777666666656679efffffeddfffffffffffffffffffffebcffffffffffffffffffffffffffffffffffffffffffff;
10'd103:marior=956'hfffffffffffffffffffffffffffffffffffffffffffedccccddbadeeeee322222221bfffffffffffffffffffecdddedea011111216fff82222213dfffffffffffffffffffffffc8888877766666655667aeffffeddfffffffffffffffffffffffbbffffffffffffffffffffffffffffffffffffffffffff;
10'd104:marior=956'hfffffffffffffffffffffffffffffffffffffffffffeddcddddbbeeeeea1222222216fffffffffffffffffffecdddeee9011112218fffa2222223cfffffffffffffffffffffffb8888877766666556667beffffedefffffffffffffffffffffffcaefffffffffffffffffffffffffffffffffffffffffff;
10'd105:marior=956'hffffffffffffffffffffffffffffffffffffffffffffddddeeeccdeeee52333223523efffffffffffffffffffcddddee7011112214fff61222122bfffffffffffffffffffffffc8888877766665556668cefffedeffffffffffffffffffffffffcaefffffffffffffffffffffffffffffffffffffffffff;
10'd106:marior=956'hffffffffffffffffffffffffffffffffffffffffffffdddeefeccddeec3233322cfb2bfffffffffffffffffffcddddde701111222159612221112afffffffffffffffffffffffd8888877666654556669ceefeedeeeeeefffffffffffffffffffcadfffffffffffffffffffffffffffffffffffffffffff;
10'd107:marior=956'hffffffffffffffffffffffffffffffffffffffffffffddefffeddddde92222224ffe27fffffffffffffffffffdddddde7011112222111222221119fffffffffffffffffffffffe8788777766645556669ceeeedddccccceffffffffffffffffffdacfffffffffffffffffffffffffffffffffffffffffff;
10'd108:marior=956'hffffffffffffffffffffffffffffffffffffffffffffeeefffeddddde61111222efb15fffffffffffffffffffdddddde7121112222221122221118ffffffffffffffffffffffff977777766554556666acdeedcccbbbccddeffffffffffffffffdacfffffffffffffffffffffffffffffffffffffffffff;
10'd109:marior=956'hffffffffffffffffffffffffffffffffffffffffffffeefffffdddddd4111111035102dffffffffffffffffffdddddde8022112222111111221118ffffffffffffffffffffffffc77776665435655566acdedccbbccccddeeffffffffffffffffcacfffffffffffffffffffffffffffffffffffffffffff;
10'd110:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffdddddd300013689aba9effffffffffffffffffeddddde9012221221111111221117fffffffffffffffffffffffff96666554356666566acdddcbcccdefffeeefffffffffffffffcacfffffffffffffffffffffffffffffffffffffffffff;
10'd111:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffdddddc46beffffffffffffffffffffffffffffedddddeb111222221111111121118ffffffffffffffffffffffffff8444433566665566acddcbccdefffffffffffffffffffffffcacfffffffffffffffffffffffffffffffffffffffffff;
10'd112:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffddddeffffffffffffffffffffffffffffffffffddddded211122211111111121109fffffffffffffffffffffffffffa66336666666566accccccceffffffffffffffffffffffffcacfffffffffffffffffffffffffffffffffffffffffff;
10'd113:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffddeffffffffffffffffffffffffffffffffffffdddddde40111221111111112101bffffffffffffffffffffffffffffe9577666666566accccccdffffffffffffffffffffffffebacfffffffffffffffffffffffffffffffffffffffffff;
10'd114:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecdddde80111121111111111003efffffffffffffffffffffffffffffc777766665566bcccccdeffffffffffffffffffffffffebadfffffffffffffffffffffffffffffffffffffffffff;
10'd115:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdddddec1111122111111111008ffffffffc6ffffffffffffffffffffe777776655566bcccccdfffffffffffffffffffffffffdbadfffffffffffffffffffffffffffffffffffffffffff;
10'd116:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdcdddde401112211111111101efffffffd417ffffffffffffffffffff977766665557bccccdefffffffffffffffffffffffffdbaefffffffffffffffffffffffffffffffffffffffffff;
10'd117:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdddddeb1111111111111000bfffffffd32329fffffffffffffffffffd77766655558cccdcdffffffffffffffffffffffffffcabefffffffffffffffffffffffffffffffffffffffffff;
10'd118:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecdddde6011111211111228fffffffc323323dfffffffffffffffffffa6666555558ccddddfffffffffffffffffffffffffebabffffffffffffffffffffffffffffffffffffffffffff;
10'd119:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdcddddd20111222102219fffffffb32333226fffffffffffffffffffd666655555accdddefffffffffffffffffffffffffdbacffffffffffffffffffffffffffffffffffffffffffff;
10'd120:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdcdddeb10111112213dfffffff9123333222cfffffffffffffffffffb66655556cccdddeffffffffffffffffffffffffecaadffffffffffffffffffffffffffffffffffffffffffff;
10'd121:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdcccdea20000114bfffffffe623333332228fffffffffffffffffffe85555559dccdedfffffffffffffffffffffffffebabeffffffffffffffffffffffffffffffffffffffffffff;
10'd122:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbcccc30159dffffffffb3233333333224efffffffffffffffffffd655547cdcddeefffffffffffffffffffffffffdaabfffffffffffffffffffffffffffffffffffffffffffff;
10'd123:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffeeeeffffffffffffc512333344333223bfffffffffffffffffffec5448dddddeffffffffffffffffffffffffffecaadfffffffffffffffffffffffffffffffffffffffffffff;
10'd124:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeffffffffffffffffffffc622333334444332229fffffffffffffffffffeeb7addddddefffffffffffffffffffffffffedbbbefffffffffffffffffffffffffffffffffffffffffffff;
10'd125:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeffffffffffffffffffa41233333344444332227fffffffffffffffffffeeeddddddddefffffffffffffffffffffffffecbacffffffffffffffffffffffffffffffffffffffffffffff;
10'd126:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeffffffffffffffc62223333334444443332226effffffffffffffffffeeeedddddddeffffffffffffffffffffffffedbbaeffffffffffffffffffffffffffffffffffffffffffffff;
10'd127:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeefffffffffffd84223333333344444443332226effffffffffffffffffeeeeeeeddddffffffffffffffffffffffffeecaabfffffffffffffffffffffffffffffffffffffffffffffff;
10'd128:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeffffffffc84223333333334444444443332226dffffffffffffffffffeeeeeeeedddffffffffffffffffffffffffedbbadfffffffffffffffffffffffffffffffffffffffffffffff;
10'd129:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeedeffeb853223333333333344444444433322227defffffffffffffffffeeeeeeeeddefffffffffffffffffffffffeebaacffffffffffffffffffffffffffffffffffffffffffffffff;
10'd130:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeedd9533223333333333334444444444333322229defffffffffffffffffeeeeeeeeeeeffffffffffffffffffffffeecbbbeffffffffffffffffffffffffffffffffffffffffffffffff;
10'd131:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeddd623333333333333344444444444333322224cdefffffffffffffffffeeeeeeeeeefffffffffffffffffffffffedbbacfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd132:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeddc623333333333333444444444433333222218ddefffffffffffffffffeeeeeeeeeeffffffffffffffffffffffeebabbefffffffffffffffffffffffffffffffffffffffffffffffff;
10'd133:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeedcc52333333333333444444444333333222223cddefffffffffffffffffeeeeeeeeeeeffffffffffffffffffffeecabadffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd134:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeddcb42333333333334444444433333322222129dddeffffffffffffffffeeeeeeeeeeeeffffffffffffffffffeeecbbacfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd135:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeedccb3233333333334444444433332222222128ccddeffffffffffffffffeeeeeeeeeeeeeffffffffffffffffeeedbbabefffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd136:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeeddcc9233333334334444444433322222222127cccddfffffffffffffffffeeeeeeeeeeedeefffffffffffffeeeecbbbaeffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd137:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeddccc623344444444444444443222222222127cccddeffffffffffffffffeeeeeeeeeeeecddeefffffffffeeeddcbbbadfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd138:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeeedddccb33444444444444444443322222211149ccccddfffffffffffffffffeeeeeeeeeeedbbcddeeeeeeeeeddddbabbbdffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd139:marior=956'hffffffffffffffffffffffffffffffffffffffffccffffffffffffffffffffffffffffffffffffffffeeeeeeddccc8244444444444444444433222211137bbcccddfffffffffffffffffeeeeeeeeeeeedbbbbcdddddddddddcbabaaefffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd140:marior=956'hffffffffffffffffffffffffffffffffffffffff69fffffffffffffffffffffffffffffffffffffffeeeeedddcccb43444444444444444443332222248bbbcccddeffffffffffffffffeeeeeeeeeeeeeda7abbbcccccccccbabbabeffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd141:marior=956'hfffffffffffffffffffffffffffffffffffffffc45ffffffffffffffffffffffffffffffffffffffeeeeedddcccc8244444444444444333333322237abbbcccddefffffffffffffffffeeeeedddeeeeeda4479abbcbbabbbbbaadffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd142:marior=956'hfffffffffffffffffffffffffffffffffffffff933bfffffffffffffffffffffffffffffffffffeeeeeeddddcccb3244444444444333333333222238abbcccddffffffffffffffffffeeeeededdeeeeeda444445555457bbaacefffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd143:marior=956'hfffffffffffffffffffffffffffffffffffffff7336ffffffffffffffffffffffffffffffffffeeeeedddddcccc61333333333333333333332222239bbcccdeffffffffffffffffffeeeeeeeddeeeeeed84444444445559bdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd144:marior=956'hfffffffffffffffffffffffffffffffffffffff6332afffffffffffffffffffffffffffffffeeeeeeddddccccc91233333333333333333322222224abccdefffffffffffffffffffeeeeeeddddeeeeeec54454444555557bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd145:marior=956'hffffffffffffffffffffffffffffffffffffffe53323efeffffffffffffffffffffffffffeeeeeedddddcccccb30232222333333333332222222226bcdeffffffffffffffffffffeeeeeeedddddeeeeea455555455555569dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd146:marior=956'hffffffffffffffffffffffffffffffffffffffd433325eeeeefffffffffffffffffffeeeeeeeedddddccccccc402222222222333333222222222229bcefffffffffffffffffffeeeeeeedddddddeeeee7455555555555568befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd147:marior=956'hffffffffffffffffffffffffffffffffffffffd4333217eeeeeeeeeeefefffeeeeeeeeeeeeedddddcccccccc601222222222222322222222222124bcceffffffffffffffffffeeeeeeeedddddddeeeec5555555555555568adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd148:marior=956'hffffffffffffffffffffffffffffffffffffffd43332228fddeeeeeeeeeeeeeeeeeeeeeedddddddcccccccc7012222222222222222222222211238ccdeeefffffffffffffffeeeeeeedddddddddeeee94555555555555568bbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd149:marior=956'hfffffffffffffffffffffffffffffffffffffff633222328eddddddeeeeeeeeeeeedddddddddcccccccccc5011222222222222222222222111227cccdeeeeefffffffffeeeeeeeeeedddddddddeeeed55555555555555569bbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd150:marior=956'hfffffffffffffffffffffffffffffffffffffff9332223327dedddddddddddddddddddddccccccccccccb5011222222222222222222221111225bcccdeeeeeeefeefeeeeeeeeeeedddddddddddeeeea45555555555555569bbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd151:marior=956'hfffffffffffffffffffffffffffffffffffffffe6222223323ceddddddddddddddccccccccccccccccca3011222222222211222222111111224bccccdeeeeeeeeeeeeeeeeeeeeeddddddddddddeeed64555555555555557abbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd152:marior=956'hffffffffffffffffffffffffffffffffffffffffe62222343217dedccccccccccccccccccccccccccc70011122222222221111111111111127cccccdeeeeeeeeeeeeeeeeeeeeedddddddddddddeef945455555555555558bbbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd153:marior=956'hffffffffffffffffffffffffffffffffffffffffff842234332118dedccccccccccccccccccccccc93011112222222222112111111111125acccccddeeeeeeeeeeeeeeeeeeedddddddddddddddeed54454555555555556abacfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd154:marior=956'hfffffffffffffffffffffffffffffffffffffffffffeb76432221026ceedccccccccccbcccccdc93001111222222222211237521111248acccccccddeeeeeeeeeeeeeeeeeedddddddddddddddeef844445555555555558bbaefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd155:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffff633221110016acdddddccccccccb85000111111222222222111269abbbbcddccccccccddddeeeeeeeeeeeeeedddddddddddddddddeefc34444554555555557ababffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd156:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffff82322111111001235778888654210011111111222222212111239aabcccccccccccccddddddeeeeeeeeeeedddddddddddddddddddeed53444445454555556abbbdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd157:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffc322211111111110000000000011111111111222222211111127bbbcccccb9cccccccdddddddeeeeeeeddddddddddddddddddddddef83444444455554556abbacfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd158:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffff82222111111112111111111111111111111111111111111127bbccccddb99bcccccddddddddddddddddddddddddddddddddddddefb3444444444445557abbabffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd159:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffd422211111111221111111111111111111111111111111126bccccddca9abbccccddddddddddddddddddddddddddddddddddddded4344444444444558abbabfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd160:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffefb2222111111122111111111111111111111111111111128ccccdddb99bccccccdddddddddddddddddddddddddddddddddddddee523333344444457abbbabefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd161:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffeefa3222111111222111111111111112321111111111126bcccdddba9bcccccccdddddddddddddddddddddddddddddddddddddee52333333444568abbbaacfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd162:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffeeeeb5222211126832211111111111259864211111237accccddca9abccccddddddddddddddddddddddddddddddddddddddddee6233344445679abbbaabdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd163:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffeeeee9521136acc921211111111116aabbcbaa9aabcdcccdcb99abcccdddddddddddddddddddddddddddddddddddddddddded63455555568bbbbbaabeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd164:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffeeeeeeedccddccccb521111111139cbbbbccccccccccccba99bcccdddddddddddddddddddddddddddddddddddddddddddddd54566555556abbaabceffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd165:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffeeeeedddddcccccccc952111137aabccccccccccccbaa99abccdddddddddddddddddddddddddddddddddddddddddddddddb545555555558bbbdefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd166:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffeeeeedddddccccccccdba9abccbba999aaaaaa999aabccdddddddddddddddddddddddddddddddddddddddddddddddccda444555545556ababfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd167:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeedddddccccccccccccccccbbbbbbbbbcccdddddddddddddddddddddddddddddddddddddddddddddddddddccdd73344444455559bbbdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd168:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeddddddcccccccccccccccccccdddddeeeeeeeeedddddddddddddddddddddddddddddddddddddddddddcccdc62344444555569bbacffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd169:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffefeeeedddddddcccccccccccccccdddeeeeeeeeeeeeedddddddddddddddddddddddddddddddddddddddddddcccdb31222222222347bbbbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd170:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffefeeedddddddddddcccdddcdcdddddeeeeeeeeeeeeddddddccccdddddddddddddddddddddddddddddddcccccd8101111211111111259ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd171:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffefeeddddddddddddddddcdcddddddeeeeeeeeedddddddcccccdddddddddddddddddddddddddddddddcccccc50011111111100001102bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd172:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffdeeedddddddddddddddddddddddddeeeedddddddcccccccdddddddddddddddddddddddddddddddcccccdb3001111111002355543100affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd173:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffddeeddddddddddddddddddddddddddddddddccccccccdddddddddddddddddddddddddddddcdccccccc7000001111013688888999854cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd174:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffdceeeddddddddddddddddddddddddddccccccccccddddddddddddddddddddddddddddddddccccccb400010111102788888889999999cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd175:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffecceedddddddddddddddddddddddddccccccdddddddddddddddddddddddddddddddddcccccccc71000100110158888898999999999aacefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd176:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdbdeeddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcccccccca30000100110378888889999999aaaabbbccefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd177:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbdeedddddddddddddddddddddddddddddddddddddddddddddddddddddddddcccccccc71000000011038888889999999aaaabbccccdddefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd178:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbdeedddddddddddddddddddddddddddddddddddddddddddddddddddddccccccbc9200000000110488888999999aaaaabcccddddeddeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd179:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbceeddddddddddddddddddddddddddddddddddddddddddddddddcccccccbbb5000000010110488889999999aaabbbccdddeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd180:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbceedddddddddddddddddddddddddddddddddddddddddddddccccccbbb8200000000011048888999999aaabbbccdddeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd181:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa439eedddddddddddddddddddddddddddddddddddddddddccccccbbba300000001101103988999999aaabbbccdddeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd182:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc633324aedddddddddddddddddddddddddddddddddddddcccccccbbba5000000000111112889999999aaabbccdddeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd183:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa323333303cedddddddddddddddddddddddddddddddddcccccccbbbb81000000000111112799999999aabbccdddeeeeeeeeeeeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd184:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd6333323300007dddddddddddddddddddddddddddddccccccccbbbbb82000000000111111069999999aaabbccddeeeeeeffeefefeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd185:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd533333410001678bdddddddddddddddddddddcdcccccccccbbbbbb94000000000001111114999999aaabbccddeeeeeeffeeefefeeeefeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd186:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc423333410003788879ddccccccccccccccccccccccccccbbbbbbb940000000001011111112899999aabbbcdddeeeeeffeefffeeefefeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd187:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa43333330000588888877addccccccccccccccccccbbbbbbbaaaa730000000000101110111179999aabbbccddeeeeeeeeeffeeefefefeeefeeeeeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd188:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa33333430001588888888778bcccbbbbbbbbbbbbbbbbbaaaaaa862000000000000011111111699aaaabbccddeeeeeeefffffefefffefefefefeeeeeefeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffffff;
10'd189:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffa43433430001689988888887778bcbbbbbbbbbbbaaaaaaaaa96300000000000101101111111389aabbbccdddeeeeffeeeeefefffefefefffefeeefefeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffff;
10'd190:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffa444434201029aa9998888888877679abbbaaaaaaaa99987410000000000000110110111111289abbbcccddeeeeeeeeefefffeeeefefefefefefefefefeefeefeeeeeeeefffffffffffffffffffffffffffffffffffffffffffffff;
10'd191:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffb44444421103abbbaaa99888888887766677898988776533100000000001010111011111111159abbcccddeeeeeeefefeeeeeefffffeffffffffffefefeefefeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffffff;
10'd192:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffc44444531103bdcccbbaaa99888888877766655544443333200100000000111111111111111148abcccddeeeeeeeeeeeeefffefeeefeffffffefffffeffefefeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffff;
10'd193:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffc44444531104eddddcccbbbaa998888887777766666555552001000101011111111111111112189bccdddeeeeeeeffeeeeeeeeffffffffeeffefefefffffffefeeffeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffffff;
10'd194:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffd54444531104deedddddcccbbbaaa99988887777766666553001010000011111111111111111159bddddeeeeeeeeeeeeeeefefeeeeeeffffffffefffffffffeffefefeeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffffff;
10'd195:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffe74444531104efeeeeeeddddccccbbbaaa9988877777666650010101111111111111111111112489cddeeeeeeeeeefeeeeeeeeeeefeffefefefeefffffeffffffffefeefeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffff;
10'd196:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffe64454531113fffeeeeeeeeeddddddcccbbbbaa99988887772011111111111111111111111122278beeeeeeeeeeeeeeeeeefeeeeeeeeeeefffffffffffffffffffeffeffefeeeeeeeeeeeefffffffffffffffffffffffffffffffffffffff;
10'd197:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffff84454531103efffeeeeeeeeeeeeeeedddddcccbbbaaa999940111111111111111111111111122589deeeeeeeeeeeeeeeeeeeeeefeffffefeffffffffffffffffffffffeffeffeeeeeeeeeeeffffffffffffffffffffffffffffffffffffff;
10'd198:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffa4555531112dfffffffeeeeeeeeeeeeeeeeeedddcccccccd81122111111111111111222222212379beeeeeeeeeeeeeeeeefeeeeeeeeeeeeeffffffeffffffefffffeffffffefefeeeeeeeeeeeeffffffffffffffffffffffffffffffffffff;
10'd199:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffb4555531111cffffffffffffffffffffffffeeeeeeffedb9521222222222222222222222222222599deeeeeeeeeeeeeeeeeeeeeeeeeeefefeffffffffffffffffffeffffffeffeffeeeeeeeeeeeefffffffffffffffffffffffffffffffffff;
10'd200:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffd65555311118ffffffffffffffffffffffffffffffdb7432222222222221112222222222222222379beeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffeeefeeeeeeeeeeeeffffffffffffffffffffffffffffffffff;
10'd201:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffff65655311118fffffffffffffffffffffffffec96431112222321248bdeedc94113222222222222599cfeeeeeeeeeeeeeeeeeeeeeeeeeeefefeffffeffffffffffffffffffffffffffefeeeeeeeeeeedfffffffffffffffffffffffffffffffff;
10'd202:marior=956'hffffffffffffffffffffffffffffffffffffffffffffff8455631111369dfffffffffffffffedba75321112223332233216dffffffffffe8222323222322379aeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefefeffffffffffffffffffffeffefffefeeeeeeeedefffffffffffffffffffffffffffffff;
10'd203:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffa56564111123333356799aa99876543222222233333333332322bffffffffffffffc42222223222599beeeeeeeeeeeeeeeeeeeeeeeeeeeeeefeefefffffffffffffffffffffffffffffffefefeeeeeeeeeeeffffffffffffffffffffffffffffff;
10'd204:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffd75551111233333332222212212222333333333333333332224efffffffffffffffff7123222222899deeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffeeffeeeeeeeeeedefffffffffffffffffffffffffffff;
10'd205:marior=956'hffffffffffffffffffffffffffffffffffffffffffffff9452111233333333333333333333333333333333332223324efffffffffffffffffff62222322399aeeeeeeeeeeeeedeeeeeeeeeeeeeeeeeeeeefeefeffffeffffffffffffffffffffffffefeeeeeeeeeeedeffffffffffffffffffffffffffff;
10'd206:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffd652111123333333333333333333333333323333333332322cffffffffffffffffffffd4123222699beeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeefefffffffffffffffffeffffffffeeeeeeeeeeeeedefffffffffffffffffffffffffff;
10'd207:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffa421111233333233233333233333332333433233333322327ffffffffffffffffffffffb122213899deeeeeeeeeeeedddeedeeeeeeeeeeeeeeeeeeeeefeeeeeeffffffffffffffffffffffffffeeeeeeeeeeeedeffffffffffffffffffffffffff;
10'd208:marior=956'hffffffffffffffffffffffffffffffffffffffffffffd631111233444333333334343343333332233333332223223dfffffffffffffffffffffee62221499aeeeeeeeeeeeeedddeeeddddedeeeeeeeeeeeeeeeeefefffeffffffffffffffffffffffffffeeeeeeeeeeeedefffffffffffffffffffffffff;
10'd209:marior=956'hffffffffffffffffffffffffffffffffffffffffffff9221112333333333333333333333333333233333322323226ffffffffffffffffffffffeea2222699aeeeeeeeeeeeeeddddeddddddeeeeeeeeeeeeeeeeeeeeeefffffefffffeffffffffffffffffffeeeeeeeeeeedeffffffffffffffffffffffff;
10'd210:marior=956'hfffffffffffffffffffffffffffffffffffffffffffc3211112333333333333333333333333333333333333332219fffffffffffffffffffffeeec2223899beeeeeeeeeeeeeddddddddddddddddeeeeeeeeeeeeeefeeeeefefffffefffffffffffffffffeeefeeeeeeeeeecffffffffffffffffffffffff;
10'd211:marior=956'hffffffffffffffffffffffffffffffffffffffffffd6211112333333233333333333333333333333333333332232afffffffffffffffffffffeedd31237a9ceeeeeeeeeeeeedddddddddddddddeeeeeeeeeeeeeeeeefefeeeeffefefefefffffffffffffffefeeeeeeeeeedcfffffffffffffffffffffff;
10'd212:marior=956'hfffffffffffffffffffffffffffffffffffffffffe73111123333333333333333333333333333333333333233332affffffffffffffffffffeeedd31223aadeeeeeeeeeeeeeeddcddddddddddddddddeeeeeeeeeeeeeeefefeeefeeeeefffffffffffffffefefeeeeeeeeeecdffffffffffffffffffffff;
10'd213:marior=956'hfffffffffffffffffffffffffffffffffffffffff9311112333333333333333332233333332333333323333233319ffffffffffffffffffffeeedc313117aeeeeeeeeeeeeeeedddcddccddddddddddeeeeeeeeeeeeeeeeeeeefeeeeeeffffffffeffffffffefeeeeeeeeeeedbefffffffffffffffffffff;
10'd214:marior=956'hffffffffffffffffffffffffffffffffffffffffb4211123343333333333333323333333333333322333323332217fffffffffffffffffffeeedcb212114beeeeeeeeeeeeeeedddccccccccddddddddddeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffeeeeeeeeeeecbfffffffffffffffffffff;
10'd215:marior=956'hfffffffffffffffffffffffffffffffffffffffc52111123333333333333333333333333333333323333233323314efffffffffffffffffeeeddca112112beeeeeeeeeeeeeeeddddcbbbbcccccddddddddddddeeeeeeeeeeeeeeefffffffffffffffffffffffeefeeeeeeeeddbdffffffffffffffffffff;
10'd216:marior=956'hffffffffffffffffffffffffffffffffffffffd6221112333333222333333333333333333333333333333233322229ffffffffffffffffeeeddcb70110218feeeeeeeeeeeeeeddddcbaabbbccccddddddddddddddeeeeeeeedefffffffffffffffffffffffffffeeeeeeeeedecbffffffffffffffffffff;
10'd217:marior=956'hfffffffffffffffffffffffffffffffffffffd63211123333333333323333333233333333333333333333322322224efffffffffffffeeeeddcba20111213dfeeeeeeeeeeeeeddddcca99aaabbcccccccccdddddddddeeeddfffffffffffffffffffffffffffffeeeeeeeeeeddbdfffffffffffffffffff;
10'd218:marior=956'hffffffffffffffffffeffffffeffffffffffd8431112233333333333333333332333333332333333233332223223227effffffffeeeeeedddcbb6011112218feeeeeeeeeeeeeddddccb989999abbbbbccccccddddddddddefffffffffffffffffffffffffffffeeeeeeeeeeeddbcfffffffffffffffffff;
10'd219:marior=956'hfffffffffffffffffffeeffeeeeeffffffed843211123332233333333323333333333333333333233333232113323218eeeeeeeeeeeedddccbb70021112212cfeeeeeeeeeeeedddddcbb8788889aaabbbbcccccdddddddffffffffffffffffffffffffffffffffeeeeeeeeedddcbeffffffffffffffffff;
10'd220:marior=956'hfffffffffffffffffffeeeeeeeeefffffed83421112333333322322333333322333333333323332333332231012323226deeeeeeeddddccbbb7001210222214feeeeeeeeeeeedddddccba857788999aaabbbcccccddcdffffffffffffffffffffffffffffffeeefeeeeeeedddccbcffffffffffffffffff;
10'd221:marior=956'hfffffffffffffffffffeeeeeeeeeffeeed9342111223333332233233333332333323333333233333333332332112322214adddddddcccbbba500122112222208feeeeeeeeeeedddddccbaa7467788999aaabbbcccccdfffffffffffffffffffffffffffffffeeeeeeeeeedddcccbbffffffffffffffffff;
10'd222:marior=956'hffffffffffffffffffffeeeeeeeeeeeed84421111233323333333333233233333333333333332233333333223210133222248abbbbbbbb9500122210112222209feeeeeeeeeeddddddccba985467778999aaabbbbbdfffffffffffffffffffffffffffffefefffeeeeeeedddccbbadfffffffffffffffff;
10'd223:marior=956'hfffffffffffffffffffffddeeeeddddc8432110122333333223333323333333333333333333333333333223233220123322222456776520012223211122222222bfeeeeeeeeeddddddccbba9854567778899aaabbdfffffffffffffffffffffffffffffffffeeeeeeeeeddddccbbacfffffffffffffffff;
10'd224:marior=956'hfffffffffffffffffffffedddddddcb833211012333333323333332333333223333333333333322333323323222220023322221111111122222222111222222211dfeeeeeeeeddddddcccba987535677778899a9dffffffffffffffffffffffffffffffffffffeeeeedddddcccbbbbfffffffffffffffff;
10'd225:marior=956'hffffffffffffffffffffffecddddd953421002333333332233232332223333323333333232232333332333323233231012332233222222232222211112212222212cfeeeeeedddddddccccba987534567777888cffffffffffffffffffffffffffffffffeeeeeeeeeeedddcccbbbbbeffffffffffffffff;
10'd226:marior=956'hffffffffffffffffffffffffdccd95542100233333333223332333333333333333332333333332332323323323333222012323222222111111111111122222222212cfeeeeedddddddccccba98765335666777cfffffffffffffffffffffffffffffffeeffeeeeeeeeddddccbbbbbbeffffffffffffffff;
10'd227:marior=956'hfffffffffffffffffffffffffecb756210023443333333233332233333332333333323333233233332332333322222232011111111100000000000111222222222211cfeeeeedddddddcccbba987653346666bffffffffffffffffffffffffffffffffffffeeeeeeeddddcccbbbbbadffffffffffffffff;
10'd228:marior=956'hfffffffffffffffffffffffffffb6521013334333332333222322232223333333333332323333233233333333323323222100000000000000000001122222223221211afeeddddddddcccccbaa8765431145bffffffffffffffffffffffffffffffffffeeeeeeeeedddddccbbbbbbadffffffffffffffff;
10'd229:marior=956'hfffffffffffffffffffffffffffd621002334333333333223333232333222323333333333333233333332322323233232231000011111212222222222222222222222217eeddddddddcccccbba986543100afffffffffffffffffffffffffffffffffffeeeeeeeeeddddccbbbbbbbadffffffffffffffff;
10'd230:marior=956'hfffffffffffffffffffffffffffd3110234333333333322222322223333232333233332323322233332332322323223223222122222222222222222222222221232221105efddddddcccccbbba987541008fffffffffffffffffffffffffffffffffeeeeeeeeeeedddddccbbabbbbadffffffffffffffff;
10'd231:marior=956'hffffffffffffffffffffffffffff700234443332333322223232233323343333233332323323233233332323333233222232232222222222222222222222222212322222118eedddddcccccbba98751007ffffffffffffffffffffffffffffffffffffeeeeeeeeddddcccbbbbabbbaeffffffffffffffff;
10'd232:marior=956'hffffffffffffffffffffffffffffe323443333332223233222323232323332323323232332333233333233333323333233222222222222222222222222222222212321222114beddccccccbbbaa851105fffffffffffffffffffffffffffffffffffeeeeeeeeeeddddcccbbbabbbbbeffffffffffffffff;
10'd233:marior=956'hffffffffffffffffffffffffffffa65544333333323222322333332323332323323333332323323333232322322333233232232222222322222222222222221222223212212114aeedcccccbba751102efffffffffffffffffffffffffffffffffeeeeeeeeeeeddddcccbbabbabbbbfffffffffffffffff;
10'd234:marior=956'hfffffffffffffffffffffffffffe7554433333333333232333223233323233332333233232333323333233332322322223223222222222322222222222222221211213212112110159bcccb96311311dfffffffffffffffffffffffffffffffffeeeeeeeeeeddddddccbbbbaabbbacfffffffffffffffff;
10'd235:marior=956'hfffffffffffffffffffffffffffa55444333333323323222322232323332333333333323232232332323323232232223322222222232222222222222222222122222212311212221101222111321519fffffffffffffffffffffffffffffffffeeeeeeeeeeedddddccbbaabbabbbadfffffffffffffffff;
10'd236:marior=956'hfffffffffffffffffffffffffff85543333333322322322223232223232323232332323333222332323223232232322323223222222232222222222222222211221112223211221111111111121146fffffffffffffffffffffffffffffffffeeeeeeeeeeeeddddcccbbaaaabbbbbefffffffffffffffff;
10'd237:marior=956'hffffffffffffffffffffffffffc6544343333222222322223332323232333233332322333222333323323222232322323223233222232222222222222221222212222121132212211111111114116effffffffffffffffffffffffffffffffefeeeeeeeeedddddcccbbaaaaabbbacffffffffffffffffff;
10'd238:marior=956'hffffffffffffffffffffffffff9554333333233223222222232323233323223333332233232332323323232232332323223233232232222222222222221222212211121211222111111111111401bfffffffffffffffffffffffffffffffffeeeeeeeeeedddddcccbbbaaaaabbbbdffffffffffffffffff;
10'd239:marior=956'hfffffffffffffffffffffffffe7544433232232222222223222222333333233332222332323323233233232222223223232222322322222222222222212212122121211112112222111111111406ffffffffffffffffffffffffffffffffeeeeeeeeeeeeddddcccbbbabababbbabfffffffffffffffffff;
10'd240:marior=956'hffffffeffffffffffffffffffc554433232222222222223232322322323223333333232322323323233232223322233232322322222222232222222222222121111212111121111222222111232dfffffffffffffffffffffffffffffffeeeeeeeeeeedddddccccbbaaaaaabbbadfffffffffffffffffff;
10'd241:marior=956'hffffffeffffffffffffffffff9554433233222222222232223232223222323233232323323333232332323323222232222323222223222222222222122121221212121111211111111111000138fffffffffffffffffffffffffffffffefeeeeeeeeeddddddccbbbaaaaaabbbbbffffffffffffffffffff;
10'd242:marior=956'hffffffefffffffffffffffffe755433333332232222322222232222332222223232332323233232332322323232232322223222222222222222222122121221211122111211111111100257889effffffffffffffffffffffffffffffffeeeeeeeeeddddddccbbbaaaaaabbbbadffffffffffffffffffff;
10'd243:marior=956'hffffffeeffffffffffffffffc65443332232322222222222223223332333323232233323333332332323323232232222323222222222222222222222121212211121111212111111105cffeeefffffffffffffffffffffffffffffffffeeeeeeeeedddddcccbbbaaaaaaabbbacfffffffffffffffffffff;
10'd244:marior=956'hffffffeeffffffffffffffffa5544332222222222222222223222323232322233222332323233232322322222232232222222223222222222222222221212211111121212111111109eeeedddffffffffffffffffffffffffffffffffeeeeeeeeedddddccccbbaaaaaaaabbbbefffffffffffffffffffff;
10'd245:marior=956'hfffffffeeeffffffffffffff8544332333222222222232223222223222222233232332323232232332322233232232222323222222222222222222221211211122111211111111108feeeeddefffffffffffffffffffffffffffffffeeeeeeeeeeddddccccbbbaaaaaaabbbadffffffffffffffffffffff;
10'd246:marior=956'hfffffffeeffffffffffffffe755343333223232222222222222223222322223232232322223232332323223232232222223222222222222222222221212211111111111111111106eeeeeeddfffffffffffffffffffffffffffffffeeeeeeeeeedddddccbbbaaaaaaaaabbabfffffffffffffffffffffff;
10'd247:marior=956'hfffffffeeffffffffffffffd65443332223222222222222222222222222223233232322223222332322323232232222322223222222222222222221212212111111111111111103ceffeeeedffffffffffffffffffffffffffffffeeeeeeeeeedddddcccbbaaaaaaaaabbbbefffffffffffffffffffffff;
10'd248:marior=956'hffffffffeefffffffffffffb65443322222222222222222222223222322232232322222232322322222232322322223222222222222222222222212122121211211111111111108eefffeeedfffffffffffffffffffffffffffffeeeeeeeeeeddddccccbbaaaaaaaaabbbadffffffffffffffffffffffff;
10'd249:marior=956'hffffffffeefffffffffffff95544333322232222222322222222222322222222222223232322322222222222322222222222222222222222222222122121111111121111111111ceeffffeedeffffffffffffffffffffffffffffeeeeeeeeedddddcccbbaaaaaaaaabbbacfffffffffffffffffffffffff;
10'd250:marior=956'hffffffffeeeffffffffffff84543323322222222222222222222223222222222222232323323222232322322222222222222222222222222222222221211111111111111111103eefffffffeefffffffffffffffffffffffffffeeeeeeeeedddddcccbbaaaaaaaaaabbabffffffffffffffffffffffffff;
10'd251:marior=956'hffffffffeeefffffffffffe75533332332222222222222222222222222222233222323323222322323223232222322222222222222222222221222212112111111111111111106eefffffffeeffffffffffffffffffffffffffefeeeeeeeedddccccbbaaaaaaaaaabbabeffffffffffffffffffffffffff;
10'd252:marior=956'hfffffffffeefffffffffffd65433333222222222222222222222222222222222223222222323322222222322222222232222322222222222222222121111111121111111111106eeffffffffeefffffffffffffffffffffffffeeeeeeeeeddddcccbbbaaaaaaaaabbbbefffffffffffffffffffffffffff;
10'd253:marior=956'hfffffffffeeeffffffffffc65443322222222222222222222222222222222222222222222223222222222222222222222222222222222222222221211111111211111111111105eefffffffffeffffffffffffffffffffffffeeeeeeeeeddddcccbbbaaaaaaaaabbbadffffffffffffffffffffffffffff;
10'd254:marior=956'hfffffffffeeeffffffffffb54433332232222222222222222222222222222222222222222222222222222222322223222222222222222221222212122111112111111111111104eeffffffffffeffffffffffffffffffffffeeeeeeeeedddddccbbbaaaaaaaaabbbadfffffffffffffffffffffffffffff;
10'd255:marior=956'hffffffffffeeefffffffff954433323222222222222222222222222222232222222222222222222222222222222222222222222222222222222221212111111111111111111101ceeffffffffffeffffffffffffffffffffeeeeeeeeedddddcccbbaaaaaaaaabbbacffffffffffffffffffffffffffffff;
10'd256:marior=956'hffffffffffeeeffffffeee954432222222222222222222222222222222222222222222222222222322222232222222222222222222222122222212122111111112111111010111aeefffffffffffeffffffffffffffffffffeeeeeeeeedddcccbbaaaaaaaaabbbacfffffffffffffffffffffffffffffff;
10'd257:marior=956'hffffffffffeeeffffeeeed7543333222222222222222222222222222222222222222222222222232222222222222222222222222222212222221212111111111111111112111106deefffffffffffefffffffffffffffffeeeeeeeeeeddddcccbabaaaaaaabbbacffffffffffffffffffffffffffffffff;
10'd258:marior=956'hfffffffffffefffeeeeeec654333332222222222222222222222222222222222222222222222232222222222222222222222222222222222121111111111112122221111111111aceeefffffffffffefffffffffffffffffeeeeeeeeddddcccbbbaaaaaaabbbacfffffffffffffffffffffffffffffffff;
10'd259:marior=956'hffffffffffffffeeeeeddb644333232222222222222222222222222222222222222222222222222222222222222222222222222222111111111111122222221121111111111114dcdeeefffffffffffeeffffffffffffeeeeeeeeeedddddccbbbaaaaaaabbbacffffffffffffffffffffffffffffffffff;
10'd260:marior=956'hfffffffffffffeeeeeddc9444333222222222222222222222222222222222222222222222222222222222222222222222211111111112212222222222121111111111111111109edbdeeeefffffffffffefffffffffffeeeeeeeeeeddddccbbbaaaaaaabbbacfffffffffffffffffffffffffffffffffff;
10'd261:marior=956'hffffffffffffeeeeddccb953333222222222222222222222222222222222222222222222222222222222222111111111112222222222222222222211121111111111111111103deecbdeeeeeffffffffffefffffffffffeeeeeeeeddddcccbbaaaaaaabbbacffffffffffffffffffffffffffffffffffff;
10'd262:marior=956'hffffffffffeeeeeddcbba875432222222222222222222222222222222222222222222222222111111111121222222223232222222222222212122111111111111111111111107eeeebbdeeeeeefffffffffeefffffefeeeeeeeeeeddddccbbbaaaaaabbbacfffffffffffffffffffffffffffffffffffff;
10'd263:marior=956'hfffffffffeeeeeddcba9996444433222211121222212111111211111111111111111211111222223334333333323222222222222222222212121111111111111111111111112ceeeeebbdeeeeeeeffffffffeeeefefefeeeeeeeeddddccbbabaaaaabbbacffffffffffffffffffffffffffffffffffffff;
10'd264:marior=956'hfffffffffeeeeddcba99d95443333333233222222222222222222222223232233223233333333333232322222232222222222222212222121211112111111111111111111106deeeeeebbddeeeeeeeefffffffeeeeeeeeeeeeeeedddcccbbbbaaaabbbacfffffffffffffffffffffffffffffffffffffff;
10'd265:marior=956'hfffffffffeedddcba99cf9444332332222222233333333222333332323333232323222232323222232222222222222222222222212222121211111111111111111111111110aeeeefeeeabcdeeeeeeeeeefffffeeeeeeeeeeeeddddcccbbbbaaaabbbacffffffffffffffffffffffffffffffffffffffff;
10'd266:marior=956'hffffffffeedddcbaa9cff9443332232222222222222222222222222232222222222222222222222222222222222222222222222121121212121211112111111111111111102deeeeeeeeebacddeeeeeeeeeeeefeeeeeeeeeeedddddcccbbbaaaabbbacfffffffffffffffffffffffffffffffffffffffff;
10'd267:marior=956'hffffffffedddcbaaabfff9543332222222222222222222222222222222222222222222222222222222222222222222222222121211212121221211111111111111111111105eeeeeeeeeeebabddddeeeeeeeeeeeeeeeeeeeeeeddddccbbbaaa9abbacffffffffffffffffffffffffffffffffffffffffff;
10'd268:marior=956'hffffffffeddcbaaaaefff8444332222222222222222222222222222222222222222222222222222222222222222222222222212122121212111111111111111111110011108eeeeeeeeefeebabcdddddeeeeeeeeeeeeeeeeedddddccbbbbaa98abbdfffffffffffffffffffffffffffffffffffffffffff;
10'd269:marior=956'hffffffffedcbaaaaeffff854333222222222222222222222222222222222222222222222222222222222222222222222222212121111111111111111111111111222221101beeeeeffefeefecaabcddddddddddeeeeeeeeeeeedcccbbbaaa889abbefffffffffffffffffffffffffffffffffffffffffff;
10'd270:marior=956'hfffffffffcbaaa9dfffff844333222222222222222222222222222222222222222222222222222222222222222221222222111211111111111111111112222222111421103deeeefefffffeffcaabccdddddddddddeeeeeeeeeeeddcbba9889aabbbfffffffffffffffffffffffffffffffffffffffffff;
10'd271:marior=956'hfffffffffcbaa9bffffff833332222222222222222222222222222222222222222222222222222222222222221212121111111111111111121222222211111111111411105eeeeeeffffffffffdaaabcccddddddddddddeeeeeeeeeeeeeeeedcbbbbdffffffffffffffffffffffffffffffffffffffffff;
10'd272:marior=956'hfffffffffeaa9afffffffa52332222222222222222222222222222222222222221222222222222122121211111111111111111212222222221111111111111111112411107eeeeeffffffffffffea9aabbccccccccccddddddeeeeeeeeeeeeeeeccbbffffffffffffffffffffffffffffffffffffffffff;
10'd273:marior=956'hffffffffffca9dfffffffa65322222222222222222222222222222222222122222222111212111111111111111111122222222221111111111111111111111111113311119eeeeeffffffffffffffb9aaabbccccccccccccddddddeeeeeeeeeddccbbefffffffffffffffffffffffffffffffffffffffff;
10'd274:marior=956'hfffffffffffabffffffffb4444432221121222222222222222212121212111111111111111111111212222232222222222212111211111111111111111111111111221111beeeeefffffffffffffffd98aaaabbbbccccccccccccdddddddddddcbbbaefffffffffffffffffffffffffffffffffffffffff;
10'd275:marior=956'hfffffffffffefffffffffc5333333333322222111121221111111111111111111122222233233323232222222121222122111211121111111111111111111111111321102ceeeeefffffffffffffffffb78aaaaabbbbbbbbbbbbbbbcccccccbbbbbbbefffffffffffffffffffffffffffffffffffffffff;
10'd276:marior=956'hfffffffffffffffffffffd5433222222222322323333232332223222332323232323222222222222212222222222122111112111111111111111111111111111111311104ceeeeeffffffffffffffffffe988aaaaaaaaaaaaaaaaaaaaaaaaaaabbbbbefffffffffffffffffffffffffffffffffffffffff;
10'd277:marior=956'hfffffffffffffffffffffd5433222222222222222222232222222222222222212121212222222222222222222221122111111111111111111111111111111111111311105deeeeeffffffffffffffffffffc8789aaaaaaaaaaaaaaaaaaaaaaaabbbbbffffffffffffffffffffffffffffffffffffffffff;
10'd278:marior=956'hfffffffffffffffffffffe7433332222222222222222232222222123112222221222121222222222222122122212121112111111111111111111111111111111111311106deeeeefffffffffffffffffffeeea878999aaaaaaaaaaaaaaaaaaaabbbacffffffffffffffffffffffffffffffffffffffffff;
10'd279:marior=956'hffffffffffffffffffffff9433332222222222222222222222222122222222222222212222222212222222222121221121111111111111111111111111111111111321107deeeeeffffffffffffffffffeeeeeb977799999aaaaaaaaaaaaaaabbbbbeffffffffffffffffffffffffffffffffffffffffff;
10'd280:marior=956'hffffffffffffffffffffffa433332222222222222222123122221222122222212221212221112221222222222211122211111111111111111111111111111111111330108deeeeeffffffffffffffffffeeeeedb98777899999aaaaaaaaaaabcbbadfffffffffffffffffffffffffffffffffffffffffff;
10'd281:marior=956'hffffffffffffffffffffffb543322222222222222222133222222122222111221122121221222212111212212111112111111111111111111111111111111111111131109deeeeeeffffffffffffffffeeeeedddb98888888999999999aaabbccbcffffffffffffffffffffffffffffffffffffffffffff;
10'd282:marior=956'hffffffffffffffffffffefd543322222222222222222223222222222222121211121212121112221212121211121111121111111111111111111111111111111111123109deeeeefffffffffffffffffeeeeedddca9988888888999999aaabbbcbcffffffffffffffffffffffffffffffffffffffffffff;
10'd283:marior=956'hfffffffffffffffffffeeee74332222222222222222122312212221322121212221212111212121211111112121111111111111111111111111111111111111111111122adeeeeeeffffffffffffffffeeeeeddcca999999999999999aaaabbbcbbffffffffffffffffffffffffffffffffffffffffffff;
10'd284:marior=956'hffffffffffffffefeeeeeef94332222222222222222212322121212121212211212121111111211112211111111111111111111111111111111111111111111111111101adeeeeeefffffffffffffffeeeeeeddccbaa99999999999aaaaaabbbcbaefffffffffffffffffffffffffffffffffffffffffff;
10'd285:marior=956'hffffffffffffffeeeeeeeefb4332222222222222222222321222121221121111121211111111211111111111112111111111111111111111111111111111111111111101bdeeeeeeefffffffffffffeeeeeeeddccbaaa999999999aaaaaaabbbcbadfffffffffffffffffffffffffffffffffffffffffff;
10'd286:marior=956'hffffffffffffeeeeeeeeeeed6323222222222222222122222222111221221121111111111121122111111111111111111111111111111111111111111111111111111101bddeeeeeeffffffffffeeeeeeeeeeddccbaaaaa9999a9aaaaaaaaabbbcacfffffffffffffffffffffffffffffffffffffffffff;
10'd287:marior=956'hfffffffffeeeeeeeeeeeeeee8432222222222222121211221111211221121211111111221111111111111111111111111111111111111111111111111111111111111101bddeeeeeeffffffffeeeeeeeeeeedddccbaaaaaaaaaaaaaaaaaaaabbbcbbfffffffffffffffffffffffffffffffffffffffffff;
10'd288:marior=956'hfffffffffeeeeeeeeeeeeeeea533222222222221222121231211111221111211211121211111111111111111111111111111111111111111111111111111111111111101addeeeeeeeeefeffeeeeeeeeeeeedddcbbaaaaaaaaaaaaaaaaaaaabbbcbbfffffffffffffffffffffffffffffffffffffffffff;
10'd289:marior=956'hfffffffffeeeeeeeeeeeeeeed633322222222222222212231221122121111211111111111111211111111111111111111111111111111111111111111111111111000000addeeeeeeeeeeeeeeeeeeeeeeeeddddcbaaaaaaaaaaaaaaaaaaaaabbbcbbeffffffffffffffffffffffffffffffffffffffffff;
10'd290:marior=956'hfffffffffeeeeeeeeeeeeeeee943322222222222211221132211111122111111111111211111111111111111111111111111111111111111111111111111111110111101addeeeeeeeeeeeeeeeeeeeeeeeeddddcbaaaaaaaaaaaaaaaaaaaaaabbbbadffffffffffffffffffffffffffffffffffffffffff;
10'd291:marior=956'hfffffffffeeeeeeeeeeeeeeeec533222222222212222221321111111221111111111111111111111111111111111111111111111111111111111111111111111111111119ddeeeeeeeeeeeeeeeeeeeeeeeedddccbabaaaaaaaaaaaaaaaaaaaabbbcbcffffffffffffffffffffffffffffffffffffffffff;
10'd292:marior=956'hfffffffffeeeeeeeeeeeeeeeee743222222222211211211321112111221111111111111111111111111111111111111111111111111111111111111111111111111211119ddeeeeeeeeeeeeeeeeeeeeeeeddddccbabaaaaaaaa999999aaaaaaabbcbbffffffffffffffffffffffffffffffffffffffffff;
10'd293:marior=956'hfffffffffeeeeeeeeeeeeeeeeeb43222222222212212211231111111121111111111111111111111111111111111111111111111111111111111111111111111222221118ddeeeeeeeeeeeeeeeeeeeeeeeddddcbbabaaaaaaaa99999999aaaaaabbbbefffffffffffffffffffffffffffffffffffffffff;
10'd294:marior=956'hfffffffffeeeeeeeeeeeeeeeeed74322222222112222222131211111121111111111111111111111111111111111111111111111111111111111111111111122222222217dddeeeeeeeeeeeeeeeeeeeeeedddccbbabaaaaaaa999999999aaaaaaabcbdfffffffffffffffffffffffffffffffffffffffff;
10'd295:marior=956'hfffffffffeeeeeeeeeeeeeeeedea5332222222222222111132111111121111111111111111111111111111111111111111111111111111111111111111111222222222116cddeeeeeeeeeeeeeeeeeeeeeddddccbaabbaaaaaa9999999999aaaaaabcbcfffffffffffffffffffffffffffffffffffffffff;
10'd296:marior=956'hfffffffffeeeeeeeeeeeeeeeeeed7432222222222122121132112111122111111111111111111111111111111111111111111111111111111111111111212222222221214cddeeeeeeeeeeeeeeeeeeeeddddccbbaabbaaaaaa9999999999aaaaaaabbbfffffffffffffffffffffffffffffffffffffffff;
10'd297:marior=956'hfffffffffeeeeeeeeeeeeeeeeedea433222222222211112123111111112111111111111111111111111111111111111111111111111111111111111122222222222212114bddeeeeeeeeeeeeeeeeeeeeddddccbbaabbaaaaa999999999999aaaaaabcbdffffffffffffffffffffffffffffffffffffffff;
10'd298:marior=956'hfffffffffeeeeeeeeeeeeeeeedddd643222222222122112113211111112111111111111111111111111111111111111111111111111111111111111222222222222221112addeeeeeeeeeeeeeeeeeeedddddccbaaabbaaaaa99998899999999aaaaabccffffffffffffffffffffffffffffffffffffffff;
10'd299:marior=956'hffffffffffeeeeeeeeeeeeeeeedddb443222222222111211122121111122111111111111111111111111111111111111111111111111111111111222222222222222222129dddeeeeeeeeeeeeeeeeeeddddccbbaaabaaaaaa999988899999999aaaabcbefffffffffffffffffffffffffffffffffffffff;
10'd300:marior=956'hffffffffffeeeeeeeeeeeeeeeddddd743222222122222211122111111112111111111111111111111111111111111111111111111111111111112222222222222222121117dddeeeeeeeeeeeeeeeeeeddddccbaaaabbaaaaa999888888999999aaaaabbcfffffffffffffffffffffffffffffffffffffff;
10'd301:marior=956'hffffffffffeeeeeeeeeeeeeeeeddddb54222222221111211114222222213111111111111111111111111111111111111111111111111111111222222222222222222221215cddeeeeeeeeeeeeeeeeeddddccbbaaaabaaaaaa9998888888889999aaaabcbdffffffffffffffffffffffffffffffffffffff;
10'd302:marior=956'hffffffffffeeeeeeeeeeeeeeeeddddd94322222222211122112312212112211111111111111111111111111111111111111111111111111112222222222222222222222114cdddeeeeeeeeeeeeeeedddddcbbaaaaabaaaaa99998888888888999aaaabbcbffffffffffffffffffffffffffffffffffffff;
10'd303:marior=956'hffffffffffedeeeeeeeeeeeeeddddddc6432222211211111111311111111211111111111111111111111111111111111111111111111111122222222222322222222222112bdddeeeeeeeeeeeeeeeddddccbaaaaaabaaaaa999888888888889999aaaabbbdfffffffffffffffffffffffffffffffffffff;
10'd304:marior=956'hfffffffffffeeeeeeeeeeeeeeeddddddb5423222221121111112211111112211111111111111111111111111111111111111111111111122222222222222232222222212119cddeeeeeeeeeeeeedddddccbaaaaaaaaaaaa99999a98777888889999aaabbbbfffffffffffffffffffffffffffffffffffff;
10'd305:marior=956'hfffffffffffedeeeeeeeeeeeeedddddcc8532222222211111111311111111311111111111111111111111111111111111111111111111222222222222222222222222221216cdddeeeeeeeeeeeeddddccbbaaaaaaaaaa999999ab98777788889999aaaabbbcffffffffffffffffffffffffffffffffffff;
10'd306:marior=956'hfffffffffffedeeeeeeeeeeeeddddddccb653332222111111111231121111221111111111111111111111111111111111111111111112222222222222222222222222222114cddeeeeeeeeeeeeddddccbbaaaaaaaaaa9999999ab97666778888999aaaaabbbefffffffffffffffffffffffffffffffffff;
10'd307:marior=956'hfffffffffffeddeeeeeeeeeeeeddddcccc954323222212211111142111111121111111111111111111111111111111111111111111222222222232222232222222222222112bcddeeeeeeeeeeddddccbbaaaaaaaaaa99999999bac98898778889999aaaabbbbfffffffffffffffffffffffffffffffffff;
10'd308:marior=956'hffffffffffeedddeeeeeeeeeedddddccccb544333222222111121231111111221111111111111111111111111111111111111111112222222222223222222222222222212119cddeeeeeeeedddddccbaaaaaaaaaaa998888989abefffffea7888999aaaaabbbcffffffffffffffffffffffffffffffffff;
10'd309:marior=956'hfffffffeeeeedddeeeeeeeeeddddddcccbb744433222222212212122111111021111111111111111111111111111111111111111122222222222232222222222222222122116cdddeeeeeeeddddccbaaaaaaaaaaa9988888889cfffffffffc889aa99aaaaabbbdfffffffffffffffffffffffffffffffff;
10'd310:marior=956'hffffffffeeedccddeeeeeeeeddddddcccbb943333333222222211214211111113111111111111111111111111111111111112111222222222222322322222222222222221213bcddeeeeeeddddccbaaaaaaaaaaa98887778889efffffffeeeb899aaaaaaaabbbbfffffffffffffffffffffffffffffffff;
10'd311:marior=956'hfffffeeeeeddeeeddeeeeeeeedddddcccbba543333333222222111114111111122111111111111111111111111111111111111122222222222222222222222222222222121129cddddeeeddddcccbaaaaaaaaaa99877677787cffffffffeeec99aaaba9aaaabbbcffffffffffffffffffffffffffffffff;
10'd312:marior=956'hfffffeeeddeffffdddeeeeedddddddcccbba543333333333222222211411111113111111111111111111111111111111111111222222222222222222322222322222221221116cddddddddddccbbaaaaaaaaaa998766666778effffffffeedcbcccccb9aaaaabbbefffffffffffffffffffffffffffffff;
10'd313:marior=956'hfffffeeeefffffffdddeeeeddddddcccbbaa633222333333322222221131112121411111111111111111111111111111122212222222222222322222322222222222222222113bcdddddddddccbbaaaaaaaa9988765555667bffffffffeedcbceeeedca9aaaabbadfffffffffffffffffffffffffffffff;
10'd314:marior=956'hfffffeeeffffffffeddeeeeddddddccbbaaa7332223333322222222221231212111411111111111111111111111111111211122222222222222232232222222222222222212118cddddddddcccbaaaaaaa998887655555668dfffffeeeeddbaceeedcba99aaaabbbfffffffffffffffffffffffffffffff;
10'd315:marior=956'hfffffeeffffffffffeeeeeddddddcccbba997333222222222222212112122112111121111111111111111111111111112212122222222222222222222222222222222212221114ccddddddcccbaaaaaaaa877666544445569fffffeeeeddcaaadddcaa9999aaabbbeffffffffffffffffffffffffffffff;
10'd316:marior=956'hfffffeeeeeffffffffeeeeddddddccbaa98763332222222222212221112112211111221111111111111111111111111121112222222222222222222232222222222222222211118cddddddccbaaaaaaaaa96555664334567cffffeeeeddcbaa8acbaaa98999aabbbeffffffffffffffffffffffffffffff;
10'd317:marior=956'hfffffddeeeefefffffeeeedddddccbaa987774332222212211211111111111211111112111111111111111111111211221222222222222222222222222322222222222222121113bcddddcccbbbbbbbaaaa8677887446668dffeeeeeddcbaaa89aaaa988999abbbbfffffffffffffffffffffffffffffff;
10'd318:marior=956'hfffffeddeeeeeeeeeefeeeddddccbaa98877642332221221111111111111111111111112111111111111111112112112211122222222222222222222232222322222222222111116cddddddddddeeeedcbaa778887667769eeefeeeddccbaa99999aa8899aabbbadfffffffffffffffffffffffffffffff;
10'd319:marior=956'hffffffdcddeeeeeeeeeeeddddccba9988777653232221211111111111111111111111111111111111101112112112211222222222222222222222222222222222222222222121111addddddddeeeeeeeedb977888677887beeeeeedddcbaaa9999aaaabbbbbbaacffffffffffffffffffffffffffffffff;
10'd320:marior=956'hfffffffccdddeeeeeeddddddccba988887766533332221111111111111000000111111111111111111110111112122112222212222222222222222223222222222222222212111115cdddddeeeeeeeeedcddca88777888aeeeeeedddcbaaaa9999aabbbaaaabcefffffffffffffffffffffffffffffffff;
10'd321:marior=956'hfffffffebccdddddddddcccbba988888777666333222221111111111111100000000111111111111111111111121221122222222222222222222222222223222222222222222111119cddddeeeeeeeeedeffffeb766789efeeeeeddccbaaa9999aabbabccdeffffffffffffffffffffffffffffffffffff;
10'd322:marior=956'hffffffffeabbcccccccbbaa999988888777777432222221111111111111111000000000000100101010101112112222121122222222222222222222222222222222222222211121113bcddddeeeeeeeeffffffffdbefffeeeeeeddccbaaaa999aaabbbeffffffffffffffffffffffffffffffffffffffff;
10'd323:marior=956'hfffffffffeaaabbbbbaa9999998888887888885333222221111111111111111001000000000000000010011111122221211222222222222222222222322222222222222222212111116ccdddeeeeeeeffffffffefffffffffedddccbaaaa9999aa9aadfffffffffffffffffffffffffffffffffffffffff;
10'd324:marior=956'hffffffffffeba9a9999999998888888888888863332222221111111111111101010000000000000000000011121222212222122222222222222222222222222222222222222221211118ccdddeeeeeeffffffffefffffffffeedccbaaaa999aaa999aefffffffffffffffffffffffffffffffffffffffff;
10'd325:marior=956'hffffffffffffcaa99999999899999888888889733222222121111111111111110100000000000000000000011112222122222222222222222222222222222222222222222212111111119ccdddeeeeeffffffffffffffffffeeebbaaaaa999aa98999adffffffffffffffffffffffffffffffffffffffff;
10'd326:marior=956'hfffffffffffffdbaaa9999aaaabaa998999aab943322222211111111111111110100000000000000000000001121222122221222222222222222222222222222222222222222211111103acddddeeeeefffffffffffffffffeeeca99aa9999a988999aadfffffffffffffffffffffffffffffffffffffff;
10'd327:marior=956'hfffffffffffffffdbabbbbbbbbaaaabbbbbbbba533232222221111111111111110101011000000000000000001122221222212222222222222222222222222222222222222222121111103bccdddeeeeeeffffffffffffffeeeeda99a989999889999aaadffffffffffffffffffffffffffffffffffffff;
10'd328:marior=956'hfffffffffffffffffecbbaabbbcdeecbaaaabbc6332322112112111111111111111100000000000000000000011222222222222222222222222222222222222222222222222212121111104acccdddeeeeeeeffffffffeeeeeddca9a989998889999aaaabdfffffffffffffffffffffffffffffffffffff;
10'd329:marior=956'hfffffffffffffffffffffeeeffffffffeeeefff73322222221211111111111111101100000000000000000000012222222222222222222222222322222222222222222222221221111111105abcccdddeeeeeeeeeeeeeeeeedddcb99899878889999aaaaabdffffffffffffffffffffffffffffffffffff;
10'd330:marior=956'hfffffffffffffffffffffffffffffffffffffff8333222222221111111111111111110000000000000000000000122222222222222222222222222222222222222222222222221212111110039abccddddeeeeeeeeeeeedddcccba88987788888999aaaaabbefffffffffffffffffffffffffffffffffff;
10'd331:marior=956'hfffffffffffffffffffffffffffffffffffffff943222222221121211111111111111000100000000000000000012222222222222222222222222222222222222222222222222221111111100179abcccddddddddddddddccbbaa988777788889999aaaaabbbfffffffffffffffffffffffffffffffffff;
10'd332:marior=956'hfffffffffffffffffffffffffffffffffffffffb433222222212121111111111111110000000000000000000000012222222222222222222222222222222222222222222222222221211111100049aabcccddddddddccccbbaaaa766777888889999aaaaabbaeffffffffffffffffffffffffffffffffff;
10'd333:marior=956'hfffffffffffffffffffffffffffffffffffffffc532222222222211111111111111111100000100000000000000002222222222222222222222222222222222222222222222222212111211100000599abbcccccccbbbaaa99aa7667777788888999aaaaabbadffffffffffffffffffffffffffffffffff;
10'd334:marior=956'hfffffffffffffffffffffffffffffffffffffffd533222222222121111111111111111100000000000000000000001222222222222222222222222222222222222222222222222222111111110000016999aaaaaaaa999999a966666677778888999aaaaabbacffffffffffffffffffffffffffffffffff;
10'd335:marior=956'hfffffffffffffffffffffffffffffffffffffffe5332222222222111211121111111110000000000000000000000001222222222222222222222222222232222222222222222222222121111110000002599999999999999aaa987766677778888999aaaaabacffffffffffffffffffffffffffffffffff;
10'd336:marior=956'hffffffffffffffffffffffffffffffffffffffff7332222222221122111112111111110000000000000000000000001222222222222222222222222222222222222222222222222221211111110000000013688988999aabbbbbbba977667777888999aaaabacffffffffffffffffffffffffffffffffff;
10'd337:marior=956'hffffffffffffffffffffffffffffffffffffffff833222222222122111111111111101101000000000000000000000132222222222222222222222222222323222222222222222222211111111101000110001125abbbbbbaabcdcbbaa87777778889999abbacffffffffffffffffffffffffffffffffff;
10'd338:marior=956'hffffffffffffffffffffffffffffffffffffffff9333222222212211112111111111110001000000000000000000001322222222222222222222222222222222222222222222222222121111111100001111111139bbaaabcdfffffedbaaa9877888899aabbadffffffffffffffffffffffffffffffffff;
10'd339:marior=956'hffffffffffffffffffffffffffffffffffffffffa332222222222212211111111111111000100000000000000000001312222222222222222222222222222222222222222222222222212111111110001111111237aceeffffffffffffedbbbaaa99aaabbbabfffffffffffffffffffffffffffffffffff;
10'd340:marior=956'hffffffffffffffffffffffffffffffffffffffffb333222222222221212111211111111100000000000000000000000202222222222222222222222222222232222222222222222222222111111111101111111225acfffffffffffffffffecbbbbbbbbbaacffffffffffffffffffffffffffffffffffff;
10'd341:marior=956'hffffffffffffffffffffffffffffffffffffffffc3332222222222121211111111111111101010000000000000000003012222222222222222222222222222222222222222222222122212111111110111111112248bffffffffffffffffffffedcbbbbbcefffffffffffffffffffffffffffffffffffff;
10'd342:marior=956'hffffffffffffffffffffffffffffffffffffffffd4332222222222212222211111111111110000000000000000000002102222222222222222222222222222222222232222222222212121111111111100111111237bdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd343:marior=956'hffffffffffffffffffffffffffffffffffffffffe5322222222222222222111111121111111000000000000000000002101222222222222222222222222222222222222222222222222222112111111111111111235acffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd344:marior=956'hfffffffffffffffffffffffffffffffffffffffff53322222222222222221221112111111111000000000000000000022002222222222222222222222222222222222232222222222222121211111111111111122349bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd345:marior=956'hfffffffffffffffffffffffffffffffffffffffff73322222222222221111111111111111111100000000000000000022001222222222222222222222222222222222222222222222222212111112111111111122348befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd346:marior=956'hfffffffffffffffffffffffffffffffffffffffff83322222222122212221211111111111111110000000000000000022001222222222222222222222222222222222222222222222222221211112111111111122236acfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd347:marior=956'hfffffffffffffffffffffffffffffffffffffffff933222222222222222221111111111111111110000000000000000120111222221222222222222222222222222222222222222222222212221211121111111222359bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd348:marior=956'hfffffffffffffffffffffffffffffffffffffffffa43322222222212222222111211111111111111000000000000000120101222222222222222222222222222222222222222222222222221212111121111111122348beffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd349:marior=956'hfffffffffffffffffffffffffffffffffffffffffb43222222222222121221112111111111111111100000000000000120111122222222222222222222222222222222222222222222222222212121221121111122347adffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd350:marior=956'hfffffffffffffffffffffffffffffffffffffffffc43322222222221222221121111111111111111101000000000000130011122222222222222222222222222222223222222222222222212122212111112111112235acffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd351:marior=956'hfffffffffffffffffffffffffffffffffffffffffd533222222222222222121111211111111111111100000000000001200011222222222222222222222222222222222222222222222222222222121211121111123348befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd352:marior=956'hfffffffffffffffffffffffffffffffffffffffffe533222222222222221211112111111111111111110000000000000201111122222222222222222222222222222222222222222222222222121212111112111122247bdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd353:marior=956'hffffffffffffffffffffffffffffffffffffffffff633222222222222222211222111111111111111111000000000000300111122222222222222222222222222222222222222222222222221222112211111211112236acfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd354:marior=956'hffffffffffffffffffffffffffffffffffffffffff7332222222222212221211111111111111111111111000000000002110111122222222222222222222222222222222222222222222222222221112121111112122349bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd355:marior=956'hffffffffffffffffffffffffffffffffffffffffff8332222222222222222111111211111111111111111000000000002101111122222222222222222222222222222222222222222222222222212111211121221122348beffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd356:marior=956'hffffffffffffffffffffffffffffffffffffffffff9323222222222212222211111111111111111111111110000000002101111222222222222222222222222222222222222222222222222222121211111111111122336acffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd357:marior=956'hffffffffffffffffffffffffffffffffffffffffffa3322222222122212121111111111111111111111111100000000021010111222222222222222222222222222222222222222222222222222222111211122122222359bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd358:marior=956'hffffffffffffffffffffffffffffffffffffffffffb4332222222222211222121112111111111111111111110000000031001111222222222222222222222222222222222222222222222222222222212111112222222348befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd359:marior=956'hffffffffffffffffffffffffffffffffffffffffffc4222222222222222221211122111111111111111111111000000021000011222222222222222222222222222222222232223222222222222212121212121122222236adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd360:marior=956'hffffffffffffffffffffffffffffffffffffffffffd43322222222222221221212111111111111111111111110000000220111112222222222222222222222222222222222222222222222222222222121212221222222349cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd361:marior=956'hffffffffffffffffffffffffffffffffffffffffffd53322222222212212222112111121111111111111111111000000220111112222222222222222222222222222222232222222222222222222222221212121122222347beffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd362:marior=956'hffffffffffffffffffffffffffffffffffffffffffe53322222222222221211121111111111111111111111111100000220111111222222222222222222222222222232222222222222222222222221212121211222222345adffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd363:marior=956'hfffffffffffffffffffffffffffffffffffffffffff632222222222121222212121111111111111111111111111100001201111122322222222222222222222222222222222223222322222222222221221222112222232349cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd364:marior=956'hfffffffffffffffffffffffffffffffffffffffffff733222222222222112222111111111111111111111111111100001201011122322222222222222222222222222222222222222222222222222221212122212222223337befffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd365:marior=956'hfffffffffffffffffffffffffffffffffffffffffff833222222222222222221221111111111111111111111111110001201111122332222222222222222222222222322222222222222222222221212121211121212222335acfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd366:marior=956'hfffffffffffffffffffffffffffffffffffffffffff9333222222222221222221211111111111111111111111111110012011111222422222222222222222222222222222222222222222222222222222211111211222222348bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd367:marior=956'hfffffffffffffffffffffffffffffffffffffffffffa333222222222122212111111112111111111111111111111110012001111112441222222222222222222222222222222222222222222222222212121212111221222236aeffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd368:marior=956'hfffffffffffffffffffffffffffffffffffffffffffa3332222222222222222121111211111111111111111111111110120011111234722222222222222222222222222222222222222222222222222222122211121212222349cffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd369:marior=956'hfffffffffffffffffffffffffffffffffffffffffffb3322222222222222121222111111111111111111111111111110020111112224842222222222222222222222222222222222222222222222222212121212122222223347befffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd370:marior=956'hfffffffffffffffffffffffffffffffffffffffffffc4332222222222221121221112112111111111111111111111111021011111223872222222222222222222222222222322222222222222222222222212212112111222336adfffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd371:marior=956'hfffffffffffffffffffffffffffffffffffffffffffd43222222222222212122121112111111111111111111111111100310111112237922222222222222222222222222222222222222222222222222212221211122222223349cfffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd372:marior=956'hfffffffffffffffffffffffffffffffffffffffffffd43222222222222222222122121111111111111111111111111110311111112236b42223222222222222222222222222223222222222222222222222212211222222223337beffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd373:marior=956'hfffffffffffffffffffffffffffffffffffffffffffe43232222222222222221212212111111111111111111111111100211111111236b72223222222222222222222222222222222222222222222222222212121212122223336adffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd374:marior=956'hfffffffffffffffffffffffffffffffffffffffffffe53322222222222222112221221111111111111111111111111101310101111236b932222222222222222222222222222222222222222222222222222221112121222223348bffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd375:marior=956'hffffffffffffffffffffffffffffffffffffffffffff63322222222222221222212121121111111111111111111111110221111112236bb51223222222222222222222222222222222222222222222222222222222222222223336aefffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd376:marior=956'hffffffffffffffffffffffffffffffffffffffffffff63322222222222211111211111111211111111111111111111110210111111235ab712222222222222222222222222222222222222222222222222222121212112222233359cfffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd377:marior=956'hffffffffffffffffffffffffffffffffffffffffffff73322222222222212222122111111111111111111111111111110221110111125aba12222222222222222222222222222222223322222222222222221221212112221222347beffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd378:marior=956'hffffffffffffffffffffffffffffffffffffffffffff73322222222222222212212121111111111111111111111111111221111111224abc32222222222222222222222222222222223222222222222222221212222222222223336adffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd379:marior=956'hffffffffffffffffffffffffffffffffffffffffffff833222222222222222212122121111111111111111111111111111101110112349bd512223222222222222222222222222222222322222222222222222221212222222223349cffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd380:marior=956'hffffffffffffffffffffffffffffffffffffffffffff843222222222222122221221111121111111111111111111111102201111112249be822222222222222222222222222222322223222222222222222222221212122222223347aefffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd381:marior=956'hffffffffffffffffffffffffffffffffffffffffffff943222222222222222222221211111111111111111111111111112201111111239bdb222222222222222222222222222222232232222222222222222222222121222222232359cfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd382:marior=956'hffffffffffffffffffffffffffffffffffffffffffff943322222222222222212112111111111111111111111111111112211111112239bce322222222222222222222222222222222222322222222222222222222122212222223348bfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd383:marior=956'hffffffffffffffffffffffffffffffffffffffffffffa43222222222122222222122111111111111111111111111111101211111112238bcf612222222222222222222222222222223222222222222222222222122222122222233346adffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd384:marior=956'hffffffffffffffffffffffffffffffffffffffffffffa43322222222222222221221111111111111111111111111111101201110111237bcf8122222222222222222222222222222222222222222223222222222212222222222233459cffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd385:marior=956'hffffffffffffffffffffffffffffffffffffffffffffa43322222222222222222221211112111111111111111111111102201111112237bbfb222222222222222222222222222222222322223222222222222222212221222222223447befffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd386:marior=956'hffffffffffffffffffffffffffffffffffffffffffffb43222222222222222222212122111111111111111111111111111211110111236abfe3222222222222222222222222223223233222232222222222222222221222222222233459cfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd387:marior=956'hffffffffffffffffffffffffffffffffffffffffffffb44322222222222222222221111111111111111111111111111112211111111236abff6122222222222222222222222222222222232322222222222222222222212222222223449bfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd388:marior=956'hffffffffffffffffffffffffffffffffffffffffffffb43322222222222222222212212111111111111111111111111112200100112236abef9122222222222222222222222222222222322322222222222222222222222122222223347adffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd389:marior=956'hffffffffffffffffffffffffffffffffffffffffffffb433222222222222222222212212111111111111111111111111022111111122359befd2222222222222222222222222222222232232232232222222222222222222222222333459cffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd390:marior=956'hffffffffffffffffffffffffffffffffffffffffffffa433222222222222222222222111111111111111111111111111122011111112349beff3122222222222222222222222222222232222232232222222222222222122222222233358befffffffffffffffffffffffffffffffffffffffffffffffff;
10'd391:marior=956'hffffffffffffffffffffffffffffffffffffffffffffa432222222222222222222222121111111111111111111111111111111101111359bdff6122222222222222222222222222222322322222322222222222222222121222222223346adfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd392:marior=956'hffffffffffffffffffffffffffffffffffffffffffff9433222222222222222222222212221111111111111111111111122111111112348bdffa2222222222222222222222222223222223223222222222222222222222222222222233358bfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd393:marior=956'hffffffffffffffffffffffffffffffffffffffffffff7433222222222222222222222222111111111111111111111111121111111112238bcffd3122222222222222222222222222222232233232222232222222222222222222222222347beffffffffffffffffffffffffffffffffffffffffffffffff;
10'd394:marior=956'hffffffffffffffffffffffffffffffffffffffffffff6332222222222222222222222221111111111111111111111111022011011122347bcfff6122222222222222222222222222222332232232232232222222222222212222222233345acffffffffffffffffffffffffffffffffffffffffffffffff;
10'd395:marior=956'hfffffffffffffffffffffffffffffffffffffffffffd5432222222222222222222222221111111111111111111111111121110111111236abfff91222222222222222222222222223223223322322222222222222222222222222222233348befffffffffffffffffffffffffffffffffffffffffffffff;
10'd396:marior=956'hfffffffffffffffffffffffffffffffffffffffffffb3323222222222222222222222211211111111111111111111111021111111112236abfffc2222222222222222222222222222222223223222222222222222222222222122222223347adfffffffffffffffffffffffffffffffffffffffffffffff;
10'd397:marior=956'hfffffffffffffffffffffffffffffffffffffffffff85443322222222222222222222221111111111111111111111111121111111112235abefff51222222221222222222222222222322322332233233222223222222222222222222333458cfffffffffffffffffffffffffffffffffffffffffffffff;
10'd398:marior=956'hffffffffffffffffffffffffffffffffffffffffffb533333333222222332222222222222211111111111111111111111211111111222359befff91222222222222222222222222222222222322222222232222222222222222222222233346aeffffffffffffffffffffffffffffffffffffffffffffff;
10'd399:marior=956'hfffffffffffffffffffffffffffffffffffffffffc5443332222223333322222222222211211111111111111111111111211111111112359bdfffd22222222222222222222222222232222223223223223322222222222222222222222233359cffffffffffffffffffffffffffffffffffffffffffffff;
10'd400:marior=956'hffffffffffffffffffffffffffffffffffffffffb44333333222222232222222222222211111111111111111111111111311111111122348bdffff41222222222222222222222222222222232233223222322222232222222222222222233347befffffffffffffffffffffffffffffffffffffffffffff;
10'd401:marior=956'hfffffffffffffffffffffffffffffffffffffffb443333233232223322233322222222221112111111111111111111111211111111122347bcffff81222222212222222222222222322322332332233223322322222222222222222222233445adfffffffffffffffffffffffffffffffffffffffffffff;
10'd402:marior=956'hffffffffffffffffffffffffffffffffffffffe5332332322222222333222332222222211211111111111111111111111211111111122347bcffffc22222222222222222222222222222223222222332232223222222222222222212222323448bfffffffffffffffffffffffffffffffffffffffffffff;
10'd403:marior=956'hffffffffffffffffffffffffffffffffffffff83333322222232222222222222222222221111111111111111111111112210111111212335abfffff51222222222222222222222222222223223222332332233222222222222222222222222346aeffffffffffffffffffffffffffffffffffffffffffff;
10'd404:marior=956'hfffffffffffffffffffffffffffffffffffffc43323322222222333332222212222222222111111111111111111111112211111111122235abeffff812222222222222222222222222222222322232223322222222222322222222222222233359cffffffffffffffffffffffffffffffffffffffffffff;
10'd405:marior=956'hffffffffffffffffffffffffffffffeeeefff9322222222222233232223222222222222111111111111111111111111132111111111222349beffffb22222222222222222222222222223222322332233222322232222222222222222222233347befffffffffffffffffffffffffffffffffffffffffff;
10'd406:marior=956'hffffffffffffffffffffffffeddcbbbbbbbabb986421122222223333222222222122221111111211111111111111111111111111111122338bdfffff412222222222222222222222222222232223322332232223222222222222222222122333359dfffffffffffffffffffffffffffffffffffffffffff;
10'd407:marior=956'hfffffffffffffffffffffdcccccccccccbbbbbbaa987421222222222332322222212222221121112111111111111111131111111111122347bcfffff912222222222212222222222222222222232223222322223222322222222222222222333447bfffffffffffffffffffffffffffffffffffffffffff;
10'd408:marior=956'hffffffffffffffffffeddcccccccccccccbbbbbaaa99986211222222333223222222122222112111111111111111111121111111111122336acfffffc22222222222222222222222222222222222232223322222222222222222222222222233346adffffffffffffffffffffffffffffffffffffffffff;
10'd409:marior=956'hfffffffffffffffffddddddddddcdccccccbbbbbaaa99999741122222222222222222122112211211111111111111112311111111111222359bffffff422222222222222222222222222222232223222222223222222222222222222222222233448cffffffffffffffffffffffffffffffffffffffffff;
10'd410:marior=956'hfffffffffffffffdddddddddddddccccccccbbbbbbaaa999997411222222222222222111211121111111111111111112211111111111222349befffff822222222222222222222222222222232232222222332223222232222222222222222333446aefffffffffffffffffffffffffffffffffffffffff;
10'd411:marior=956'hfffffffffffffedddddddddddddccccccccccbbbbbaaaa99999973112222222222222111122111111111111111111112111111111121223337adfffffc222222222222222222222222222222222322332233222332232222222222222233233334569cfffffffffffffffffffffffffffffffffffffffff;
10'd412:marior=956'hffffffffffffedddddddddddddddddccccccccbbbbbaaaa9999999731112222222222111112211111111111111111113211111111111122346acffffff522222222222222222222222222222222222222332223322322222222222222222212335557beffffffffffffffffffffffffffffffffffffffff;
10'd413:marior=956'hfffffffffffedddddddddddddddddddccccccccbbbbbaaaa999999996212222222221211111221111111111111111112111111111111222335abffffff8123222222222222222222222222223222222232223322222222222222222222222222223469dffffffffffffffffffffffffffffffffffffffff;
10'd414:marior=956'hffffffffffddddddddddddddddddddddccccccccbbbbbaaaaa99999898401112222221111111121111111111111111121111111111111123349befffffc322222222222222222222222222232223223322233222223223222222222222122122122247bffffffffffffffffffffffffffffffffffffffff;
10'd415:marior=956'hfffffffffddddddddddddddddddddddddcccccccbbbbbbaaaaa9999999983111122112211121111211111111111111121111111111121223348beffffff5222222222222222222222222222222322332233222223223322222222222122112112122237dfffffffffffffffffffffffffffffffffffffff;
10'd416:marior=956'hffffffffdddddddddddddddddddddddcccccccccbbbbbbaaaa99999999899611111221112111111111111111111111221111111111111122336bdffffff82223322222222222222222222222232223233222222323322322322222122111211111222247fffffffffffffffffffffffffffffffffffffff;
10'd417:marior=956'hfffffffedddddddddddddddddddddddccccccccbbbbbbbaaaaaa9999999889830111122111211111111211111111111111111111111111223358cffffffc2223222222222222222222222223322322332222222332332222222222221121111111121224affffffffffffffffffffffffffffffffffffff;
10'd418:marior=956'hffffffecddddddddddddddddddddddddccccccccbbbbbaaaaaaaa999999898996111111112111111111121111111111111111111111121222335afffffff42232322222222212222222222222232232222233332332222222211111122111112111121234bfffffffffffffffffffffffffffffffffffff;
10'd419:marior=956'hffffffdddddddddddddddddddddddddddccccccccbbbbaaaaaaaaa999999999997301111111111111111112111111112111111111111111222347cffffff622332222222222222222222222222232232232333223222222212221111111111111111112236dffffffffffffffffffffffffffffffffffff;
10'd420:marior=956'hfffffddddddddddddddddddddddddddccccccccccbbbbbbaaaaaa99999999988899501111111111111111111111111221111111111111122223459efffff9222322222222222222222222222222233233233233222222211211111111100000001111111139efffffffffffffffffffffffffffffffffff;
10'd421:marior=956'hfffffcddddddddddddddddddddddddddcccccccccbbbbbbaaaaaa99999989988888983011111111111111111112111221111111111111222222348bfffffc3223222222222222222222222222223223333232222222211211111100002456899aaaabbbbbaabdefffffffffffffffffffffffffffffffff;
10'd422:marior=956'hffffdcdddddddddddddddddddddddddddccccccccbbbbbbbaaaa999999988988888888511111111111111111111112121111111111221222122337bdffffd3223222222222222222222222222222223332222222222221111000135899aaaaaaaaabbbbbbbbbbbbbcefffffffffffffffffffffffffffff;
10'd423:marior=956'hfffeccddddddddddddddddddddddddddccccccccbbbbbbbaaaaa999999999988888888972011111111111111111111232212111211111111122237bcffffe42223222222222222222222222332222332332322222111110001579aaaaaaaaaabbbbbbbbbbbbbbbbbbabcdffffffffffffffffffffffffff;
10'd424:marior=956'hfffdcccddddddddddddddddddddddddddcccccccbbbbbbaaaaaaa99999998988888888889500111111111111111111132111111111111111112249bbfffff622232222222222222222222332222222332222222111100037abaaaaaaaaabbbbbbbbbbccbbbbbbbbbbbbbabcffffffffffffffffffffffff;
10'd425:marior=956'hfffccccddddddddddddddddddddddddddcccccccbbbbbaaaaaaa99999999989888988888897301111111111111111113211111111111111111235abbfffff5222322222222222222222222223222223222222111001379aaaaaaaaabbbbbbbbbbbbccccccccccbbbbbbbbbabdffffffffffffffffffffff;
10'd426:marior=956'hffebccccccddddddddddddddddddddddddcccccbbbbbbaaaaaaa99999999998888988888888861011111111111111112211111111111111111237bbcfffff5232232222222222222223322322222222222211100169aaaaaaabbbbbbbbbccccccccccccccccccccccbbbbbbbabdffffffffffffffffffff;
10'd427:marior=956'hffdccccccccdcddddddddddddddddddddcdccccccbbaaaaaaaaaa999999889888888888888888840011111111111111121111111111111111225abadffffc3222332222222222222342222222222222222110048baaaaaaaabbbbbbbbbbccccccccccccccccccccccbbbbbbbbbaceffffffffffffffffff;
10'd428:marior=956'hffccccccccccccddddddddddddddddddddcccccccbbbaaaaaaaa999999889988888888888888888730011111111111122111101111111111224abbbeffff922222322222222222243222222222222212110039aaaaaaaaabbbbbbbbccccccccccccccccccccccccccccbbbbbbbbabefffffffffffffffff;
10'd429:marior=956'hfecbcccccccccccdddddddcddddddddddcccccccbbbbaaaaaaaa999999888888888888888888888896300010010111111011000010111111357abacfffff4223224222222222234222222222222211110039baaaaaaabbbbbbbbbbbcccccccccccccccccccccccccccccccbbbbbbaadffffffffffffffff;
10'd430:marior=956'hfdbbbccccccccccccccccddcdddddddcccccccccbbbbaaaaaaa99999998888888888888888888888889741001011000210101101111112456779bbfffffd22222233222222223322222222222221111038baaaaaaaabbbbbbbbbcccccccccccccccccccccccccccccccccccbbbbbbaabfffffffffffffff;
10'd431:marior=956'hfcbbcccccccccccccccccddddddddcccccccccccbbbbaaaaaaa99999988888888888888888888888888887432110000201111111122456666678acfffffa222222432222222322222222222221111017bbaaaaaaabbbbbbbbbccccccccccccccccddddddddddccccccccccccbbbbbbaabffffffffffffff;
10'd432:marior=956'hfcbbbbbbcccccccccccccccccccccccccccccccbbbbaaaaaaaa99999888888888888888888888788888888875443333212222334556666666678abfffff623223322222222322222222222221111039baaaaabbbbbbbbbbbbbcccccccccccccddddddddddddddccccccccccccbbbbbbaabeffffffffffff;
10'd433:marior=956'hfbbbbbbbbbbcbccccccccccccccccccccccbcccbbbaaaaaaaaa99999888888888888888888888888888888878765555555555555555566666677aaefff93322222332222332222222222221111017baabaaabbbbbbbbbbbbcccccccccddddccdddddddddddddddcccccccccccccbbbbaaaaefffffffffff;
10'd434:marior=956'hebbbbbbbbbbbbccccccccccccccccccccccbbbbbbbaaaaaaaa999999888888888888888888888888888788877877655555555555555666666677aadfff5243232232222232222222222121111039baaaaaabbbbbbbbbbbccccccccccdddddddddddddddddddddddccccccccccccbbbbaaaabfffffffffff;
10'd435:marior=956'heabbbbbbbcbbbbcbbcbcccccccccccccccccbbbbbbaaaaaa999999988888888887888888888888888887877777778765555555555666666666779bcffc32233333322222222222222111111005bbaaaaaabbbbbbbbbbccccccccccddddddddddddddddddddddddddccccccccccccbbbbaaaabffffffffff;
10'd436:marior=956'heaabbbbbbbbbbbbbbbbbbccbccccccbcbbbcbbbbbbbaaaaa99999999888888888888888778778787777877777777777766555555666666666667abcff93232222222223222222222111111018baaaaaaaabbbbbbbbccccccccccccddddddddddddddddddddddddddccccccccccccbbbbaaaaabfffffffff;
10'd437:marior=956'hdaabbbbbbbbbbbbbbbbbbbbbbccbbbbbbbbbbbbbbaaaaaaa99999998888888888887887777777777777777777777777777666555566666666667abcff7333222232223222222222111111039aaaaabbbbbbbbbbbbbccccccccccccddddddddddddddddddddddddddccccccccccccbbbbaaaaaacffffffff;
10'd438:marior=956'hdaabbabbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbabaaaaa999999988888888888887787777787777777777777777777777776665666666666668abcff83333222222222222221211111105aaaabbbabbbbbbbbbbbbcccccccccccdddddddddddddddddddddddddddccccccccccccbbbbbaaaa9adfffffff;
10'd439:marior=956'hdaaaaaaabbbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaaaaaaa999999888888888888887777777777777777777777777777777766666666666666668aacffa433222342222222212111111017aaaaabbbabbbbbbbbbbbcbcccccccccdddddddddddddddddddddddddddcccccccccccccbbbbbaaaa99aeffffff;
10'd440:marior=956'hdaaaaaaabbbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaaaaaa9999998888887888888877777777777777777777777776776766666666666666666668badffc53333333222222211211210128aaaaabaabbbbbbbbbbbbbccccccccccccddddddddddddddddddddddddddcccccccccccccbbbbbaaaa99acffffff;
10'd441:marior=956'heaaaaaaaaabaaabbbaabbbbbbbbbbbbbaaaaaaaaaaaaaa9999988888888888877777777777777777777677776766766666666666666666666679badfff6333324322221221111111149aaaaabbabbbbbbbbbbbbbbccccccccccccdddddddddddddddddddddddddccccccccccccccbbbbbbaaa999aefffff;
10'd442:marior=956'hea9aaaaaaaaaaabaabaaaaaaabbbaabbaaaaaaaaaaaa99999998898888888887777777777777777777667666666666666666666655655666667abaefffb4333233112221111110125aaaaaaaabbbbbbbbbbbbbbbbcccccccccccddddddddddddddddddddddddcdcdccccccccccccbbbbbaaaa9999bfffff;
10'd443:marior=956'hfa99aaaaaaaaaaaaabbaaaaaaaaaaaaaaaaaaaaaaa9999999998898888888777777777777777677776776666666666666666655565656666668bbbfffff733223412221121111236aaaaaaaaababbbbbbbbbbbbcbcccccccccddddddddddddddddddddddddddccccccccccccccbbbbbbbaaaa9999adffff;
10'd444:marior=956'hfb999aaaaaaaaaaaaabaaaaaaaaaaaaaaaaa9aaaa99999999998888888888877777777777776677666666666666666666665555555556666669bacffffff6333232122111122348aaaaaaaaaabbbbbbbbbbbbbbbbcccccccccddddddddddddddddddddddddddccccccccccccbbbbbbbbbaaaa9999abffff;
10'd445:marior=956'hfb9999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa99999999999888888888888877777667776667666666666666665555665555555555566667abbdffffffd63223311112233359aaaaaaaaaaaaaabbbbbbbbbbbbcccccccccddddddddddddddddddddddddccdccccccccccccbbbbbbbbbaaaa99989bdfff;
10'd446:marior=956'hfc98999999a99aaaaaaaaaaaaaaaaaaaaaaa9aa999999999999888888888877777777677666666666666665666665555665565555555556669bbbeffffffd865424423444446aaaaaaaaaaaaaaaabbbbbbbbbbbbccccccccdddddddddddddddddddddddddccccccccccccbbbbbbbbbbbbaaa999989acfff;
10'd447:marior=956'hfe9889999999999a9aaaaaaaaaaaaaaaaaaa99999999999999888888888877777776666666666666666666556665555556555555555555667abacfffffffd97666665555568aaaaaaaaaaaaaaaaabaabbbbbbbbbccccccccdddddddddddddddddddccddccccccccccccccbbbbbbbbbbbaaaa9999889bfff;
10'd448:marior=956'hffa888889999999999999999aaaa9aaaa9a99999999999999888888888777777777666666666666666666655666656555555555555555557abbbefffffffda97666666668aaaaaaaaaaaaaaaaaaababbbbbbbbbbcccccccddddddddddddddddddcccccccccccccccccbbcbbbbbbbbbbaaaa99999889adff;
10'd449:marior=956'hffc8888888898899999999999aa99a999999999999999888888888888777777777776666666666666666665555665555555555555555557abbadffffffffd99987666689aaaaaaaaaaaaaaaaaaabbbbbbbbbbbbcccccccdddddddddddddddddccccccccccccccccccbbbbbbbbbbbbbaaaaa99999889acff;
10'd450:marior=956'hfff87888888888998899999999999999999999999999988888888888777777777666666666666666666666666555555555555555555668abbabfffffffffd999aaa99aaaaaaaaaaaaaaaaaaaaababbbbbbbbcccccccccccccdcddddddddddccccccccccccccccccccbbbbbbbbbbbbbaaaa999998888abef;
10'd451:marior=956'hfffb7778888888888889899999999999999999999988888888888887777777776666666666666666666666666555555555555555567889abbbffffffffffe9999aaaaa9aaaaaaaaaaaaaaaaaaaaaaaabbbbbbbcbccccccccccccddcddcdcccccccccccccccccccccbbbbbbbbbbabbaaaaa999998888abdf;
10'd452:marior=956'hffff9777778888888888888899999988888998888888888888888777777777766666666666666666666666566555555555555677888999abacffffffffffe99999999999aaaaaaaaaaaaaaaaaaaaaaabbbbbbbcbccccccccccddddccccccccccccccccccccccccbbbbbbbbbbbaaaaaaaaaa999988889bcf;
10'd453:marior=956'hffffe87777777778888888888888888888888888888888888777777777777776666666666666666666666555655555566677888899999aabacfffffffffffa99999999a9aaaaaaaaaaaaaaaaaaaabbbbbbbbbbbcbbbccccccccddcccdcccccccccccccccbbcbbbbbbbbbbbbbaaaaaaaaaa9998888889acf;
10'd454:marior=956'hfffffd767777777777778888888888888888888888777777777777777766666666666666666666566556555556667777888889999999aaabacfffffffffffb89999999999aaaaaaaaaaaaaaaaaaaaabbbbbbbbbbccbccccccccccccccccccccccccccccbbbbbbbbbbbbbbbaaaaaaaaaa999998888888abf;
10'd455:marior=956'hffffffd76667777777777788888877788878777777777777777667666666666666666666666665565565556677788888889999999999aaabacfffffffffffc99999999999999aaaaaaaaaaaaaaaaaabbbbbbbbbbbccccccccccccccccccccccccbcccbbbbbbbbbbbbbbbaaaaaaaaaaaa999988888788abe;
10'd456:marior=956'hfffffffe96666777777777777787777777777777777777777766666666666666555655656665655555667878888889999999999999aaabbbacfffffffffffe999999999999999aaaaaaaaaaaaaabbbbaaabbbbbbbbccccccccccccccccccccccbbbbbbbbbbbbbbbbbbaaaaaaaaaaa999999988888778abe;
10'd457:marior=956'hffffffffb976666666777777777777777777766666666666666666666666555555555555655665566788877889999999999999aaaabbbbbabfffffffffffffa8999999999999aaaaaaaaaaaaaaabbbaabbbbbbbbbbbbbbbccccccbbcccccbccbbbbbbbbbbbbbbbabbbaaaaaaaaaa9999999888887778abe;
10'd458:marior=956'hffffffffdcb87665666666677777776777776776666666666666666655555555555555555555567788877789999999999999aaabbbbaaabdffffffffffffffc8899989999999a9aaaaaaaaaaaaabaaaabbbbbbbbbbbbbcccbbbbbbccccbbbbbbbbbbbbbbbbbbaaaaaaaaaaaaaa999999998888887778abd;
10'd459:marior=956'hffffffffeeeeca9766556666666666666666666666666666666555555555555555555555556788889998778999999aaaaabbbbbbaaabdefffffffffffffffff98889889999999999aaaaaaaaaaaaaaaaabbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbabbbbaaaaaaaaaa999999999988888877778bbd;
10'd460:marior=956'hffffffffeeeeeeeca987655555666666666666666665555555555555555555555555555677888999abbaa989aaaaabbbbbbaaabbcdfffffffffffffffffffffb8888888999999999aa99aaaaaaaaaaaaabbbabbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbaaabaaaaaaaaaaa99999999999888888777778bbd;
10'd461:marior=956'hffffffffeeeeeeeffedca9765555555555555555555555555555555555555555555567888889999abbbabaabbbbbbaaaaabcdefffffffffffffffffffffffffe9888888999999999999aaaaaaaaaaaaaaabaaabaabbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaaaaaaaaaaa9999999999988888887777779bbe;
10'd462:marior=956'hffffffffeeefffffffffffedcb9876555555445555555555555555555554555667888899999999abbbadfedbaabbbcdeffffffffffffffffffffffffffffffffc888888898999999999aaaaaaaaaaaaaaaaaaaaaaaabbabbbbbbbbbbbbbbbbbbbaaaaaaaaaaaaaaa99a9999999999888888877777789bbe;
10'd463:marior=956'hfffffffffeeffffffffffffffeeedcba98877666555555555555555556677888889999999999aabbbbdffffffefffffffffffffffffffffffffffffffffffffffa7888888899999999a9aaaaaaaaaaaaaaaaaaaaaaaaaabbbbbbaababaabaaaaaaaaaaaaaaaaaa999999999999998888887777777789bbe;
10'd464:marior=956'hffffffffffcdffffffffffffffeeeeeeeedccba998888888888888888899999999999999999abbbabeffffffffffffffffffffffffffffffffffffffffffffffff878888888889999999999aaaaaaaaaaaaaaaaaaaaaaaaaabaaaaaaaaaaaaaaaaaaaaaaaaaa999a99a999999999888888777777778abbf;
10'd465:marior=956'hffffffffffebbceffffffffffffffeeeeeeeeeeeddcbba99999999999999999999999999aabbbbabffffffffffffffffffffffffffffffffffffffffffffffffffe87888888888999999999aaaaaaaaaaaaaaaaaaaaaaaaaaabaaaaaaaaaaaaaaaaaaaaaa9999a99999999999999888887777777778abbf;
10'd466:marior=956'hffffffffffffcbabcdefffffffffffeeeeeeeeeeeddddddccbaa99999999999999999aaabbbbabdffffffffffffffffffffffffffffffffffffffffffffffffffffa87777888888999999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa9aaa9aa9aaaa99999999999999988888887777777778abcf;
10'd467:marior=956'hffffffffffffffdbaabbceeffffffffeeeeeeeeeeedddddddddccbaa999999999aaaaabbbbaacffffffffffffffffffffffffffffffffffffffffffffffffffffffda887777888889999999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa999a99999999999988888888888777777777779bacf;
10'd468:marior=956'hfffffffffffffffffdbaaaabcdeeeeffeeeeeeeeeeddddddddccccccbaaaaaaaaabbbbbaabdffffffffffffffffffffffffffffffffffffffffffffffffffffffffddb98877788888999999999aaaaa9aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa999999999999999998888888888877777777777779badf;
10'd469:marior=956'hffffffffffffffffffffdcbaaaabbbcccdddeeeededdddddddcccccbbaaaaaabbbbbaabceffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddeda98877888889999999999999aa99aaaaaaaaaaaaaaaaaaaaaaaaa999a999999999999999998888888888877777777777777abbef;
10'd470:marior=956'hfffffffffffffffffffffffedcbaaaaaaaaabbbbbbbbbbbbbbaaaaaaaabbbbbaaaabdefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeddeeb9998788888899999999999a9999aaaaaaaaaaaaaaaaaaaaa9999999999999999999999898888888887777777666667778abbff;
10'd471:marior=956'hffffffffffffffffffffffffffffedccbbaaaaaaaaaaaabbbbbbbbbbbaaaabbcdeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeeeeeea99987888889999999999999aa9aaaa9aaaaa9aaaaa99aaaaaaa99999999999988888888888888877777776666666779bacff;
10'd472:marior=956'hfffffffffffffffffffffffffffffffffffeddcccbbbbbbbbbbbbbbbccddeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddeeeec99988888999999999999999aa99aa9999aaa99aa99aa9999999999999999989898888888887777777766666666677abadff;
10'd473:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcceeeeda9988888899999999999999999999999aaaa9999a999999999999999988888888888887777777776666666666678bbbfff;
10'd474:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdabdefeb9778888898889999999999999999a9aaa99aa9999999999999999998888888888888777777766666666666667abacfff;
10'd475:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffebabcefc7798788888888999999999999999999999a99999999999999988888888888887777777767766666666666668bbbdfff;
10'd476:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffebaabda79a87788888888898899999999999999999999999999998888888888888877777776666666666666666667abacffff;
10'd477:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbaabbca877788888888888899998899899988899999988888888888888877777777767666666666666666667abbbeffff;
10'd478:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbacda87777888888888888888888888888888889888888888888877777777777766666665566556666669bbacfffff;
10'd479:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedddb877778778888888888888888888888888888888888877777777776666666666655555555566668bbabffffff;
10'd480:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeddc9766777777777887888888888888888888878777777777777776666666655555555555666669bbbbeffffff;
10'd481:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedddca8666777777788777777788888878777777777777777666666666665555555555555555669bbbadfffffff;
10'd482:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeddddb9766667777777777777777777777777777776666666666666555555555555555555568abbbadffffffff;
10'd483:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddeeedb9766666777777777777777777767776666666666666665555555555555555555679bbbabdfffffffff;
10'd484:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffddeeeedb9765666666666666666666666666666666666665555555555555555555566789abbabeffffffffff;
10'd485:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedeeeeeeeca8765556666666666666666666666555555555555555555555555566789999abbaefffffffffff;
10'd486:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedeeeeeeeedca87665555556666666656565555555555555555555555556678889999aaabbaefffffffffff;
10'd487:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedeeeeeeeeeedcb987665555555555555555555555555555555566778888999999aaaaabbaefffffffffff;
10'd488:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeceeeeeeeeeeeeedcba9877766555555555555555666777788889999999999aaaaaaaabbaefffffffffff;
10'd489:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecdeeeeeeeeeeeeeeeddca99888888888888888888889999999999999aaaaaaaaaaabbbbffffffffffff;
10'd490:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbbdeeeeeeeeeeeeeeeeeeddcba99888899999999999999999aaaaaaaaaaaaaaaabbbacffffffffffff;
10'd491:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdabdeeeeeeeeeeeeeeeeeeeeeeeddcbaa99999aaaaaaaaaaaaaaaaaaaaaaaaabbbabfffffffffffff;
10'd492:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbbcdeeeeeeeeeeeeeeeeeeeeeeeeeddccbbaaaaaaaaaaaaaaaaaaaaaaabbbbabffffffffffffff;
10'd493:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecaabcdefeeeeeeeeeeeeeeeeeeeeeeddddddcbbaaaaaaaaaaaaaaabbbbaabdfffffffffffffff;
10'd494:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdbaaabcdeeeeeeeeeeeeeeeeeeddddddddddddccbaaaaaaabbbbbaaabdfffffffffffffffff;
10'd495:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbaaabbbccdeeeeeeeeeeeddddddddcccbbbaaaabbbbbbaaabcdffffffffffffffffffff;
10'd496:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedbaaaaaabbbbbcbbcbbbbbbbbaaaaaaabbbbbaaaaabcdefffffffffffffffffffffff;
10'd497:marior=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdcbbaaaaaaaaababbabbbbbaaaaaaaabbccdeffffffffffffffffffffffffffff;
10'd498:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeddcbbbbbbbbbbbbbbcccddeefffffffffffffffffffffffffffffffffff;
10'd499:marior=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
	endcase

	case((y_cnt-move_y))
10'd0:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeedba98777666789abcdefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd1:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec9754332222222222222222334579befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd2:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc964222222222222222222222222222222346adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd3:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda6322222222222221121111111111222222222222236adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd4:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffea63222222222222211111111111111111111112222222222359dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd5:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7322222222222221211111111111111111111111111111222222226bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd6:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb532222222222222222111111111111111111111111111111112222222227cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd7:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffb6322222222222222222212111111111111111111111111111111111222222235bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd8:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffd73222222222222222222212111111111111111111111111111111111111122222224afffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd9:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffff832222222222122222221222221111111111111111111111111111111111111122222224afffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd10:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffc532222222221111111112221111111111111111111111111111111111111111111112222224bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd11:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffff8322222221100135677642001111111111111111111111111111111111111111111111122222225cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd12:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffe722222221025aefffffffffeb520111111111111111111111111111111111111111111111122222227dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd13:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffd6322222103aeffdccccccdcdfffe920111111111111111111111111111111111111111111111122222239ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd14:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffd422222103cffdcdeffffffbeeddefff80011111111111111111111111110010111111111111111122222225cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd15:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffb42222212affddfffffffffa39fffdceffe30111111111111111111101111100000101111111111111112222238fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd16:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffc43222113efddffffffffffd544effffddefe50111111111111111110110100000000001011111111111112222225cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd17:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffd43222107fedefffffffffff74427fffffedeff601111111111111111111010010000000001011111111111122222239ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd18:mariog=956'hffffffffffffffffffffffffffffffffffffffffffd5222211afedffffffffffffa44344cffffffceff501111111111111111110000000000000000011111111111112222226dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd19:mariog=956'hffffffffffffffffffffffffffffffffffffffffff63222118fde5affffffffffc5443437fffffffcdfe301111111111111111000000000000000000001011111111112222224cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd20:mariog=956'hfffffffffffffffffffffffffffffffffffffffff83222108fefc439fffffffff64443343bfffffffdefc0111111111110110101000000000000000000001011111111112222239ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd21:mariog=956'hffffffffffffffffffffffffffffffffffffffffa3322107feff94539fffffffa444433333cfffffffdff60111111111111000000000000000000000000010111111111112222226effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd22:mariog=956'hfffffffffffffffffffffffffffffffffffffffd5222113feefd544538fffffd54444333336fffffffeefd10111101011111100000000000000000000000000111111111112222225efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd23:mariog=956'hfffffffffffffffffffffffffffffffffffffff6322211bfeffb4445446ffff744444333333afffffffdef601111111101000000000000000000000000000000011111111111222224bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd24:mariog=956'hffffffffffffffffffffffffffffffffffffff93222107fefff843444447dfb4444433333334dffffffeefb100101001001000000000000000000000000000000101111111111222233afffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd25:mariog=956'hfffffffffffffffffffffffffffffffffffffd4322112defffe6434444447e744444323334437fffffffefe30111111000000000000000000000000000000000000011111111112222339ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd26:mariog=956'hfffffffffffffffffffffffffffffffffffff73221108fefffc44334444445444443333333333affffffeee600000000010000000000000000000000000000000000001111111112222338fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd27:mariog=956'hffffffffffffffffffffffffffffffffffffa4222111deffff843334444444444432c923333334cfffffeef9000000000000000000000000000000000000000000000011111111112222337ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd28:mariog=956'hffffffffffffffffffffffffffffffffffff63221105fefffe543334444444444435fd333333335ffffffefb0000000000000000000000000000000000000000000000001111111111222337fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd29:mariog=956'hfffffffffffffffffffffffffffffffffffa3322111aeffffc44333234444444433cff7233333336fffffeec10000000000000000000000000000000000000000000000000111111112222336ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd30:mariog=956'hfffffffffffffffffffffffffffffffffff63221113eeffffa44332853444444326fffd233333333cffffdec200000000000000000000000000000000000000000000000001111111112222336effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd31:mariog=956'hffffffffffffffffffffffffffffffffffb33221105feffff844332cf534444432bffff5233333335dfffeed2000000000000000000000000000000000000000000000000001111111112222337ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd32:mariog=956'hffffffffffffffffffffffffffffffffff632211109fffffe633333dfe52444434fffffb3333333336fffefd20000000000000000000000000000000000000000000000000010111111111222336fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd33:mariog=956'hfffffffffffffffffffffffffffffffffb43221110bfffffd533333dfff5334429ffffff6233333333afffec200000000000000000000000000000000000000000000000000001111111111222337ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd34:mariog=956'hfffffffffffffffffffffffffffffffff832211111ceffffa433324efffd42433effffffb2333333333bffeb1000000000000000000000000000000000000000000000000000000011111112222338fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd35:mariog=956'hffffffffffffffffffffffffffffffffe532211102deffff7333324effffe5228ffffffff62333333335deda00000000000000000000000000000000000000000000000000000000111111111222338ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd36:mariog=956'hffffffffffffffffffffffffffffffffa332211102eefffe6333325fffffff42dffffffffc22333333327fe800000000000000000000000000000000000000000000000000000000011111111222334afffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd37:mariog=956'hffffffffffffffffffffffffffffffff7332111102defffc4433326fffffffe9ffffffffff7233333322bfd7000000000000000000000000000000000000000000000000000000000011111111222334cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd38:mariog=956'hfffffffffffffffffffffffffffffffd5322111102defffb4333327fffffffffffffffffffd32333331afdc40000000000000000000000000000000000000000000000000000000000011111111122235cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd39:mariog=956'hfffffffffffffffffffffffffffffffb3322111101defffa4433327fffffffffffffffffeff92333326eeda100000000000000000000000000000000000000000000000000000000000011111111222336effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd40:mariog=956'hfffffffffffffffffffffffffffffff93322111101beeff73333328ffffffffffffffffeeefe423324deed70000000000000000000000000000000000000000000000000000000000000011111111222337ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd41:mariog=956'hffffffffffffffffffffffffffffffe632211111109efff74333328fffffffffffeeeeeeeeeeb2223cdeeb300000000000000000000000000000000000000000000000000000000000000101111111222338fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd42:mariog=956'hffffffffffffffffffffffffffffffd532211111106fefe53333329ffffffffeffeeeeeeeeede511acdfd9100000000000000000000000000000000000000000000000000000000000000001111111122234affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd43:mariog=956'hffffffffffffffffffffffffffffffb432211111003eefc4333332afffffffeeeeeeeeeeedddda16dcfdb50000000000000000000000000000000000000000000000000000000000000000000111111122234cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd44:mariog=956'hffffffffffffffffffffffffffffff9332211110100afec4333332affeeeeeeeeeeeeedddddcdd9bbeec8100000000000000000000000000000000000000000000000000000000000000000001111111122336dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd45:mariog=956'hffffffffffffffffffffffffffffff73322111110005eeb3433332bfeeeeeeeeeeeddddddddcdddcdeca40000000000000000000000000000000000000000000000000000000000000000000001111111122337efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd46:mariog=956'hffffffffffffffffffffffffffffff63222111100000cfc3233332bfeeeeeeeddddddccccddeeeeedca6000000000000000000000000000000000000000000000000000000000000000000000011111111222349fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd47:mariog=956'hfffffffffffffffffffffffffffffe532211111100004efe732332aeeeeddddddcddeeeeeeddddccca71000000000000000000000000000000000000000000000000000000000000000000000001111111122234bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd48:mariog=956'hfffffffffffffffffffffffffffffd4322111110000009eeeb5222aedddddcccdeedddcccba9865433211100000000000000000000000000000000000000000000000000000000000000000000001111111122236dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd49:mariog=956'hfffffffffffffffffffffffffffffc4322111100000001bffed9309ddddccdefecccba8643322333332211111000000000000000000000000000000000000000000000000000000000000000000011111111122238effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd50:mariog=956'hfffffffffffffffffffffffffffffb43221111100000001ceeddd89cccdeeedcb974333333333333333222111111010000000000000000000000000000000000000000000000000000000000000011111111112224affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd51:mariog=956'hfffffffffffffffffffffffffffffa432211111000000002beedccccceedca8543344444433333223322221111111111111110000000000000000000000000000000000000000000000000000000001111111112236dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd52:mariog=956'hfffffffffffffffffffffffffffff93322111110000000001adeecbdfdb75434444433333333333322222221111111111111111111000000000000000000000000000000000000000000000000000001111111112238dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd53:mariog=956'hfffffffffffffffffffffffffffff7332211110000000000006bdefd9643444444444333332222222222222221111111111111111111110000000000000000000000000000000000000000000000000111111111222458effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd54:mariog=956'hfffffffffffffffffffffffffffff733221111100000000000038a74334444333322222211122111111111111111111111111111111111111000000000000000000000000000000000000000000000001111111112234358effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd55:mariog=956'hfffffffffffffffffffffffffffff7332111111000000000000123333333222222221111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111112244334afffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd56:mariog=956'hfffffffffffffffffffffffffffff633221111000000000012343322222222111111000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000001011111111123433336cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd57:mariog=956'hfffffffffffffffffffffffffffff6332211110000000013333222211100000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000111111111223333334bffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd58:mariog=956'hffffffffffffffffffffffffffffe633221111100001233222211110000000000000000000100110000000000000000000000000000001111112111111110000000000000000000000000000000000000001111111112333333349fffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd59:mariog=956'hffffffffffffffffffffffffffffe6332211100012332221110000000000000011111111111111111111111111111100000000000000000001111111111111000000000000000000000000000000000000011111111112322233348ffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd60:mariog=956'hffffffffffffffffffffffffffffe63322110123322110000000000000111111111111111111111111111111111111111111110000000000000011111111111100000000000000000000000000000000000101111111122222233338fffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd61:mariog=956'hffffffffffffffffffffffffffffe633211233311100000000000011111111111111111111111111111111111111010000000111111000000000000011211111110000000000000000000000000000000000111111111122222223338ffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd62:mariog=956'hfffffffffffffffffffffffffffff6322333210000000000011111111111111111111111111111111111111111100100000000001111111000000000001111111111000000000000000000000000000000000111111111122222223349fffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd63:mariog=956'hfffffffffffffffffffffffffffff6344311000000000111111111111111111111111111111111111111111111100000000000000000001111000000000001111111110000000000000000000000000000000011111111111122222335cffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd64:mariog=956'hfffffffffffffffffffffffffffff73210000000011111111111111111111111111111111111111111111111100000000000000000000011101111000000000111111110000000000000000000000000000001011111111111122222337dfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd65:mariog=956'hfffffffffffffffffffffffffffc6100000000111111111111111111111111111111111111111111112223333444444331000000000000000000011110000000011211110000000000000000000000000000000011111111111112222349effffffffffffffffffffffffffffffffffffffffffffffffff;
10'd66:mariog=956'hffffffffffffffffffffffffff820000000111121111111111111101111111111111111111122344455555555555554310000000000000000122111111110000001111111100000000000000000000000000000001111111111111222236bffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd67:mariog=956'hffffffffffffffffffffffffb30000000111222111111111111010111111111111111123445555555555555555555430000000000000000000144443211111110000011111100000000000000000000000000001010011111111111222348efffffffffffffffffffffffffffffffffffffffffffffffff;
10'd68:mariog=956'hfffffffffffffffffffffff8100000011222111111111111111000001111111111234455555555555555555555554300000000000000000000024444444322111100011121111000000000000000000000000000001001111111111122235bfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd69:mariog=956'hfffffffffffffffffffffe600000111222211111111111111100000001111112344555555555555555556666655530000000000000000000000034454544443211110011122110000000000000000000000000000000101111111111122349dffffffffffffffffffffffffffffffffffffffffffffffff;
10'd70:mariog=956'hffffffffffffffffffffd3000000122221122111111111110000000011012345555555555555656666666666665400000000000000000000000014555555544443211101112211000000000000000000000000000001110111111111122237befffffffffffffffffffffffffffffffffffffffffffffff;
10'd71:mariog=956'hfffffffffffffffffffd30000012222112222111111111100000000011244555555555555666666666666666665100000000000000000000000003555555555444432111111121100000000000000000000000000000000011111111122235adfffffffffffffffffffffffffffffffffffffffffffffff;
10'd72:mariog=956'hffffffffffffffffffd3000011222212222111111111110000000000244555555555566666666666666666666530000000000000000000000000015555555555554443111111111100000000000000000000000000000001011111111122249bfffffffffffffffffffffffffffffffffffffffffffffff;
10'd73:mariog=956'hfffffffffffffffffd20000112221222221111111111100000000024455555555666666666666666666666666410000000000000000000000000004556665555555554431121101110000000000000000000000000000000001111111122238beffffffffffffffffffffffffffffffffffffffffffffff;
10'd74:mariog=956'hfffffffffffffffff500001122212222221111111111000000001344555555666666666666666666667776766200000000000000000000000000002566666666555555554311110000000000000000000000000000000000110111111112236adffffffffffffffffffffffffffffffffffffffffffffff;
10'd75:mariog=956'hffffffffffffffff8000111221122222212111111110000000122334555566666666666666666677777777765100000000000001233332100000000566666666666655555542100000000000000000000000000000000000001011111112235acffffffffffffffffffffffffffffffffffffffffffffff;
10'd76:mariog=956'hfffffffffffffffb2000111211222221211111111100000001100002455666666666666777777777777777764000000000012456666677665310000466676666666666666655420000000000000000000000000000000000000011111112234abffffffffffffffffffffffffffffffffffffffffffffff;
10'd77:mariog=956'hfffffffffffffff500111121122222122211111111000000100000000355666666666777777777777777777620000000014566677777777777641003677777777776777777666520000000000000000000000000000000000000111111112349befffffffffffffffffffffffffffffffffffffffffffff;
10'd78:mariog=956'hffffffffffffffd200111121122222222111111110000001000000000025666666777777777777777777777510000001366777777777777777787301677777777777777777777640000000000000000000000000000000000000001111112249bdfffffffffffffffffffffffffffffffffffffffffffff;
10'd79:mariog=956'hffffffffffffff7111111111122222222111111110000010000000000002566677777777777777777777777400000026777787888888888777777851677777777777777788887761011110000000000000000000000000000000001111112249bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd80:mariog=956'hfffffffffffffe3001111111122221211211111100000100000000000000366777777777777777777777777400000377788888888888888888887786788777777788888888888873011111110000000000000000000000000000001111112248bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd81:mariog=956'hfffffffffffffd3111111111211112112111111110001100000000000000056777777777777777777777777300004788888888888888888888888888888888888888888888888885001111111100000000000000000000000000011111112248bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd82:mariog=956'hfffffffffffffb2111111112112122111111111110002000000111110000026777777777777777777777777200047888888888888888888888888888888888888888888888888886011111111111000000000000000000000000001111112248bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd83:mariog=956'hfffffffffffffa1111111111111111111111111100012000001111111000005777777777777777888888887200378888888888888888888888888888888888888888888888999887101111111112210000000000000000000000000111112249bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd84:mariog=956'hfffffffffffffb2011111111111111111111111010022000111111111100003677777777777788888888887202688888888888888888888888888888888888888888888899999988201111111112222000000000000000000000000111112249bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd85:mariog=956'hfffffffffffffc2111111111111111111111111100031001111111111110001677777788888888888888887205888888888888888888888888888888888888888888889999999988201111111112222200000000000000000000011111112249bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd86:mariog=956'hfffffffffffffd311111111111111111111111000014001111111111111100047777888888888888888888823888888888777888778888888888888888888888888999999999999830111111111222222000000000000000110000011111235abcfffffffffffffffffffffffffffffffffffffffffffff;
10'd87:mariog=956'hffffffffffffff6111111111111111111111111000240011123445544321100378888888888888888888888479888888789abbbcba977888999999999999888888899999999999983011111111122222220000000004789abba974100111236aacfffffffffffffffffffffffffffffffffffffffffffff;
10'd88:mariog=956'hffffffffffffffa1111111111111111111111000003401114566666666542101688888888888888899999a99a9999878abcccccccccb9889aaaaaaaaaaaaaaaa999999999999999830111111111222222210000017abbbbbbbbbbcc82011237badfffffffffffffffffffffffffffffffffffffffffffff;
10'd89:mariog=956'hffffffffffffffe3111111111111111111111100004401146677777777765310588888888888999aaaaaaaaaaaa9879bccccccccccccca89aabbbbbbbbbbbbbbbaaaaaaaa9999998301111111112222222200004aaaabbbbbbbbbbbbb601238bbdfffffffffffffffffffffffffffffffffffffffffffff;
10'd90:mariog=956'hfffffffffffffffa11111111111111111111110000540136777777788887763038888888999aaaaabbbbbbbbaaa989cccdddddddddddddb8aabbbbbbbbbbbbbbbbbbbbbbaaaa999941111111111122222221006aabbbbbbbbbbbbbbbbc81249bbefffffffffffffffffffffffffffffffffffffffffffff;
10'd91:mariog=956'hffffffffffffffff81111111111111111111100000550267777778888888876327888999aaaabbbbbbbbbbbaaa989bdddddddededddedddc9abbbbbbbbbbbbbbbbbbbbbbbbaaaa994111111111112222222106abbbbbbbbbbbbbbbbbbbc924abbffffffffffffffffffffffffffffffffffffffffffffff;
10'd92:mariog=956'hfffffffffffffffff5111111111111111111100000550577777888888888888757999aaaabbbbbbbbbbbbbbaaa98bdddeeeeeeeeffeeeeedb9abbbbbbbbbbbbbbbbbbbbbbbbaaa99411111111112222222103abbbbbbbbbbbbbbbbbbbbbb95abcffffffffffffffffffffffffffffffffffffffffffffff;
10'd93:mariog=956'hffffffffffffffffff5111111111111111111100005627777888888888888888889aaaabbbbbbbbbbbbbbbbaa98acdeeeeeeeefc7422359dda9bbbbbbbbbbbbbbbbbbbbbbbbaaaa9411111111112222222128bbcbbbbbbbbbaaabbbbbbbbbaaadffffffffffffffffffffffffffffffffffffffffffffff;
10'd94:mariog=956'hfffffffffffffffffff8211111111111111111100067677888888888877888899aaaabbbbbbbbbbbbbbbbbbaa99bdeeeeeeefb4223444433bd9abbbbbbbbbbbbbbbbbbbbbbbaaaa931111111111222223215abcbbbbbbaaaaaaaaaaabbbbbbbaeffffffffffffffffffffffffffffffffffffffffffffff;
10'd95:mariog=956'hffffffffffffffffffffb4111111111111111111006777888888888769aaa9899aaaaaabbbbbbbbbbbbbbbbaa9acdeeeeeefa234566667642ac9bbbbbbcbbbbbbbbbbbbbbbbbaaa821211111112222223228bcbbbbbaaa99988899aaaababbbbfffffffffffffffffffffffffffffffffffffffffffffff;
10'd96:mariog=956'hfffffffffffffffffffffd8411111111111111110068888888888866bcccccba9aaaabbbbbbbbbbbbbbbbbbaa9bdeeeeeefa14577777787543b9abbbccbbcbbbbbbbbbbbbbbbaaa72221111122222222324abbbbbbaa988877777899aaaababbeffffffffffffffffffffffffffffffffffffffffffffff;
10'd97:mariog=956'hffffffffffffffffffffffec9742211111111111106988888888875bcccccddca9aaaabbbbbbbbbbbbbbbbba99bdeeeeeec3467887778966644aabbbbcccccbbbbbbbbbbbbbbaa951222211112222222326abbbbbaa98887777777899aaaaabbcffffffffffffffffffffffffffffffffffffffffffffff;
10'd98:mariog=956'hffffffffffffffffffffffffdbba976555567875207988888888759cccdddddeebaaaabbbbbbbbbbbbbbbbba99cdeeeeee636778888898677536abbbccccbccbbbbbbbbbbbbbaa832222221222222223328abbbbaa988888888888889aaaaaabbefffffffffffffffffffffffffffffffffffffffffffff;
10'd99:mariog=956'hffffffffffffffffffffffffffecbbbbbbbbbbbb927a9888888866ccdddddeeb988aaabbbbbbbbbbbbbbbbba9acdeeeeec3578889866778876538abbccccccbcbbbbbbbbbbbbaa622222221222222223339abbbaa98888889aaa999899aaaaabbcfffffffffffffffffffffffffffffffffffffffffffff;
10'd100:mariog=956'hfffffffffffffffffffffffffffffeccbbbbbbbbc76a9888888759dddddeeb42224aaabbbbbbbbbbbbbbbbba9adddeeef736898a7332226877746abbcccccbbcbbbbbbbbbbbbaa422222222222222223349aabaa988889aaaaaaaa9999aaaaaabbeffffffffffffffffffffffffffffffffffffffffffff;
10'd101:mariog=956'hffffffffffffffffffffffffffffffffffffffffffaa998888875bdddddea3345547aabbbbbbbbbbbbbbbbba9bdddeeee43689a733222225887659bbbccbbcbcbbbbbbbbbbbba9322222221222222223349aaaa998889aaaaaaaaaa999aaaaaabbdffffffffffffffffffffffffffffffffffffffffffff;
10'd102:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffb999888865dddddeb34677766aaabbbbbbbbbbbbccbba9bdddddec2577992229ec422788659bbbbccccbbbbbbbbbbbbbba7222222222222222223359aaaa9888aaaaaaaaaaaaa999aaaaabbcffffffffffffffffffffffffffffffffffffffffffff;
10'd103:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffc999888867edeeee4577777669aabbbbbbbbbbccbcbba9bdddddea146785117fff922598768bbbbbbbbbbbbbbbbbbbbbba7233222222222222223469aaa99889aaaaaaaaaaaaaa99aaaaabbbffffffffffffffffffffffffffffffffffffffffffff;
10'd104:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffca99999979eeeeea4787886668aabbbbbbbbbbccccbba9bddddde9156893118fffb22279857abbbbbbbbbbbbbbbbbbbbba6232222222222322223479aaa9889aaaaaaaaaaaaaaaaaaaaaabbaefffffffffffffffffffffffffffffffffffffffffff;
10'd105:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffda999aa97aeeeee66899733646aabbbbbbbbbcccccbba9bddddde8156882215fff712158877abbbbbbbbbbbbbbbbbbbbbb7232222222222211223579aaa989aaaaaaabbbabbaaaa9aaaaabbaefffffffffffffffffffffffffffffffffffffffffff;
10'd106:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffda99aaaa8bddeec5789732dfb28babbbbbbbbcccccbba9bddddde72468722226a7222149876abbbbbbbbbbbbbbbbbbbbbb8222222221222111223589aa988998999aabbbbbbbbaaaaaaaaabadfffffffffffffffffffffffffffffffffffffffffff;
10'd107:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffeaaaaaaa8cddde95887325fff35babbbbbbbcccccccba9bddddde7256872222111222239976abbbbbbbbbbbbbbbbbbbbbb9222222222222111223589aa98887777789abbbbbbbbaaaaaaaabacfffffffffffffffffffffffffffffffffffffffffff;
10'd108:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffebaabbaa9cddde74796123efc14abbbbbbbbcccccccbb9bddddde7145772222222222227876abbbbbbbbbbbbbbbbbbbbbba41222221122111222368999887666666679abbbbbbbbaaaaaaabacfffffffffffffffffffffffffffffffffffffffffff;
10'd109:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffbabbbba9ddddd65784111462129abbbbbbbcccccccbbaaddddde8146882222221122227976abbbbcbbbcbbbbbbbbbbbbbb711111111111111223689998777777777779abbbbbbbaabaaaabacfffffffffffffffffffffffffffffffffffffffffff;
10'd110:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffcbbbbbaaddddd5687235677887abbbbbbbbcccccccbbaacdddde9035783122111112227a87abbbccccccbbbbbbbbbbbbbba41111111012112223689987777789999888abbbbbbbaabaaaabacfffffffffffffffffffffffffffffffffffffffffff;
10'd111:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffcbbbbbaaddddc68bbcccccbbbbbbbbbbbbbcccccccbbaacdddddb134584122111111227987abbccccccccccccbbbbbbbbbba401110011111122368987777899aaaaa989abbbbbbaabaaaabacfffffffffffffffffffffffffffffffffffffffffff;
10'd112:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffdbbbbbaaddddcbbbbbbbbbbbbbbbbbbbbbbcccccccbbaabdddddc225697122111111128977bbcccccccccccccccbcbbbbbbba5210012221122237888778899aaaabaa99abbbbbbaabaaaabacfffffffffffffffffffffffffffffffffffffffffff;
10'd113:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffecbbbba9ccbbbbbbbbbbbbbbbbbbbbbbbbbbbcccccbbaabddddde425688121111111129a78bbccccccccccccccccbbbbbbbbaa8312222211222378887888aaaaaabba999bbbbbcbbbaaaabacfffffffffffffffffffffffffffffffffffffffffff;
10'd114:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffecbbbbabbbbbccccccccccccccbbbbbbbbbbbbbccbbbaaaccddde81457b41111111114b879bcccccccdcccbbbbbbbbbbbbbbbaa712222111122378888889aaaaabbbba99bbbbbcbbbaaaabadfffffffffffffffffffffffffffffffffffffffffff;
10'd115:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffcbbbbccccccccccccccccccccccccbbbbbbbbbbbcbbbaacccdddb2358a81111111117b98bccccccc84bbbbbbbbbbbbbbbbbbba92222211112237888888aaaaaabbbba99bbbbbcbbbaaabbadfffffffffffffffffffffffffffffffffffffffffff;
10'd116:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffcbbcccccccccccccccccccccccccccbbbbbbbbbbbbbbaabcccddd41679b511111103ba79bccbbbc9204bbbbbbbbbbbbbbbbbbba4122211112248888889aaaaabbbbbaa9bbbbbcbbbaaabbaefffffffffffffffffffffffffffffffffffffffffff;
10'd117:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffdbccccccccccccccccccccccccccccccbbbbbbbbbbbbaaacccccda1479ab5011103bba9abbbbbc911216cbbbbbbbbbbbbbbbbbb8222221112248898889aaaabbbbbbaaabbbbccbbaaaabbbefffffffffffffffffffffffffffffffffffffffffff;
10'd118:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffdcccccccccccccccccccccccccccccccccbbbbbbbbbbaaabcccccd61689ac84237bba9abbbbbb82122129bbbbbbbbbbbbbbbbbba51211111225889888aaaabbbbbbbaaabbbbcccbaaaabbbffffffffffffffffffffffffffffffffffffffffffff;
10'd119:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffecccccccccccccccccddddccccccccccccbbbbbbbbbbbaaabccccdc13689bbccccb99aaaaabc811222214bbbbbbbbbbbbbbbbbbb92111111226989989aaaabbbbbbbaaabbbcccbbaaaabacffffffffffffffffffffffffffffffffffffffffffff;
10'd120:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffdcccccccccccccccddddddddddccccccccccbbbbbbbabbaaabccccdb1269aabbba9aaaaaabb60122222218bbbbbbbbbbbbbbbbbbb6111111238889989aaabbbbbccbaabbbccccbaaaabbbdffffffffffffffffffffffffffffffffffffffffffff;
10'd121:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffdccccccccccccccdddddddddddddccccccccccbbbbbbaabbaaabccccda214678889aaaaaaba412222222215bbbbbbbbbbbbbbbbbbba311111269889989aaabbbbcccbaabbcccccbaaaabbbeffffffffffffffffffffffffffffffffffffffffffff;
10'd122:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffcccccccccccccccddddddddddddddcccccccccbbbbbbaaabaaaabbbcccc401479aaaaaabb811222222221129bbbbbbbbbbbbbbbbbab921111499989a9aaabbbbcccbaabccccccbaaaaababfffffffffffffffffffffffffffffffffffffffffffff;
10'd123:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffdcccccccccccccccddddddddddddddcccccccccbbbbbbbaaabaaaabbbbbbbabbbaaaaabb83112222222221127bbbbbbbbbbbbbbbbbbaa81115999989a9aabbbbbbcbaabccccccbbaaaabbadfffffffffffffffffffffffffffffffffffffffffffff;
10'd124:mariog=956'hffffffffffffffffffffffffffffffffffffffffffeccccccccccccccccddddddddddddddcccccccccbbbbbbbaaaaaaabbbabaaaaaaaaabbb8311222222222221215baabbbbbbbbbbbbbbbaaa846a999999aaabbbbbbbbbabcccccccbbaaaabbbefffffffffffffffffffffffffffffffffffffffffffff;
10'd125:mariog=956'hffffffffffffffffffffffffffffffffffffffffffdccccccccccccccccccddddddddddddcccccccccbbbbbbbaaaaaaabbbbabaaabaabca7211222222233322211139babbbbbbbbbbbbbbbaaaaa99999999aabbbbbbbbbbbbbcccccbbaaaabbacffffffffffffffffffffffffffffffffffffffffffffff;
10'd126:mariog=956'hffffffffffffffffffffffffffffffffffffffffffdccccccccccccccccccddddddddddddcccccccccbbbbbbbaaaaaaabbbbbbbbbbba8411122222222333322211138aaababbbbbbbbbbbbaaaaaaaa9999abbbbbbbbbbbbbbbccccbbaaa9abbaeffffffffffffffffffffffffffffffffffffffffffffff;
10'd127:mariog=956'hfffffffffffffffffffffffffffffffffffffffffecccccccccccccccccccddddddddddddccccccccbbbbbbbbaaaaaaabbbbbbbbb9521112222222233333222211137aaaabbbbbbbbbbbaaaaaaaaaaa999abbabbbbbbbbbbbbcccbbbaa9abbabfffffffffffffffffffffffffffffffffffffffffffffff;
10'd128:mariog=956'hfffffffffffffffffffffffffffffffffffffffffdcccccccccccccccccccccdddddddddcccccccccbbbbbbbaaaaaaaabbbcca85211122222222223333332222211379aaaabbbbbbbbbbbaaaaaaaaaa999abbbbbbbbbbbbbbbbcbbbaaa9abbadfffffffffffffffffffffffffffffffffffffffffffffff;
10'd129:mariog=956'hfffffffffffffffffffffffffffffffffffffffffdcccccccccccccccccccccdcdddcccccccccccccbbbbbbbaaaaa999aa852111122222222222333333322222111479aaaabbabbbbbbbaaaaaaaaaaaa99abbbbbbbbbbbbbbbbbbbaaa9abbacffffffffffffffffffffffffffffffffffffffffffffffff;
10'd130:mariog=956'hfffffffffffffffffffffffffffffffffffffffffdccccccccccccccccccccccccccccccccccccccbbbbbbbbaaaaa99521111222222222222223333333222222111588aaaaabbbbbbbbbaaaaaaaaaaaaaaabbbbbbbbbbbbbbbbbbaaa99bbbbeffffffffffffffffffffffffffffffffffffffffffffffff;
10'd131:mariog=956'hfffffffffffffffffffffffffffffffffffffffffccccccccccccccccccccccccccccccccccccccbbbbbbbbaaaaa998411222222222222222333333332222221112678aaaaaabbbbbbbbbaaaaaaaaaaaaaabbbbbbbbbbbbbbbbbaaaa9abbacfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd132:mariog=956'hffffffffffffffffffffffffffffffffffffffffeccccccccccccccccccccccccccccccccccccccbbbbbbbbaaaaa998411222222222222223333332222222111114778aaaaaabbbbbbbbbaaaaaaaaaaaaaabbbbbbbbbbbbbbbbaaaa9abbbbefffffffffffffffffffffffffffffffffffffffffffffffff;
10'd133:mariog=956'hffffffffffffffffffffffffffffffffffffffffeccccccccccccccccccccccccccccccccccccbbbbbbbbbaaaaa9998312222222222222233333322222222111126778aaaaaaabbbbabbaaaaaaaaaaaaaaaabbbbbbbbbbbbbaaaaa99bbbadffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd134:mariog=956'hffffffffffffffffffffffffffffffffffffffffecccccccccccccccccccccccccccccccccccbbbbbbbbbaaaaaa9988212222222222222333332222222211111157788aaaaabbbbaabbaaaaaaaaaaaaaaaaaaabbbbbbbaaaaaaa999bbbacfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd135:mariog=956'hfffffffffffffffffffffffffffffffffffffffffcccccbccccccccccccccccccccccccccbbbbbbbbbbbaaaaaa99987222222222222223333222222211111111477889aaaabababbabaaaaaaaaaaaaaaa9aaaaaaaaaaaaaaaaa999abbabefffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd136:mariog=956'hfffffffffffffffffffffffffffffffffffffffffccccbbbbcccccccccccccccccccccbbbbbbbbbbbbbaaaaaaa9988612222222222233333322222211111110377788aaaaababaabbaaaaaaaaaaaaabaa999aaaaaaaaaaaaa9999abbbaeffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd137:mariog=956'hfffffffffffffffffffffffffffffffffffffffffdbbbbbbbbbccbcccccccccccbbbbbbbbbbbbbbbbbaaaaaaa99988312222222222233333222211111111103777888aaaaaaabbbaaaaaaaaaaaaaaabaa88899aaaaaaaaa99999abbbadfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd138:mariog=956'hfffffffffffffffffffffffffffffffffffffffffdcbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaa999988722222333333333333322221111111015777888aaaaaaaaaaaaaaaaaaaaaaaaaabaa767889999999999889abbbbdffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd139:mariog=956'hffffffffffffffffffffffffffffffffffffffffbacbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaaa999988513223333333333333222221111101367778889aaaaaaababaaaaaaaaaaaaaaaabba7667888888888889abbbaaefffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd140:mariog=956'hffffffffffffffffffffffffffffffffffffffff57cbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaaa9999988722322333333332222222221111114677778889aaaaaaaaabaaaaaaaaaaaaaaaabbb964667777788889abbbbabeffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd141:mariog=956'hfffffffffffffffffffffffffffffffffffffffb34cbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaaaaa999988851322233332332322222222111136667778889aaaaaaaaaaaaaaaaaaaaaaaaaaabbba711356778877abbbbaadffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd142:mariog=956'hfffffffffffffffffffffffffffffffffffffff8229cbbbbbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaaaaa999998887113222232222222222222221111466777888aaaaaaaaaaaaaaaaaaaaaaaaaaaaabbba6111112222236bbaacefffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd143:mariog=956'hfffffffffffffffffffffffffffffffffffffff6225cbbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaaaaaaa999998888402222222222222222222221111256777789aaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbba41111111112239cdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd144:mariog=956'hffffffffffffffffffffffffffffffffffffffe52218cbbbbbbbbbbbbbbbbbbbabaaaaaaaaaaaaa9999999888860122222222222222222221111112677789aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbb921111111112225bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd145:mariog=956'hffffffffffffffffffffffffffffffffffffffd42212bbaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa99999998888720121212222222222222211111113779aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbb7111111111112249dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd146:mariog=956'hffffffffffffffffffffffffffffffffffffffc322214bbaaaaaaaaaaaaaaaaaaaaaaaaaaaaa999999988888830111111112222222221111111111577aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbb4111111111112237befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd147:mariog=956'hffffffffffffffffffffffffffffffffffffffc3222216baaaaaaaaaaaaaaaaaaaaaaaaa9999999999888888300111111111122222111111111112778aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbb91111111111112237adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd148:mariog=956'hffffffffffffffffffffffffffffffffffffffd32221116baaaaaaaaaaaaaaaaaaaaaa999999999888888884001211111111111111111111111115888aaaaaaaaaaaaaaaaaaaaaaaaaa9aaaaaaaabbb51111111111112237bbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd149:mariog=956'hfffffffffffffffffffffffffffffffffffffff522212216baaaaaaaaaaaaaa9999999999999888888888830011111111111111111111111111037888aaaaaaaaaaaaaaaaaaaaaaaa9a9aaaaaaabbba11111111111111238bbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd150:mariog=956'hfffffffffffffffffffffffffffffffffffffff9222112225aa9999999999999999999999988888888888300111111111111111111111111110278889aaaaaaaaaaaaaaaaaaaaaa9999999aaaaabbb601111111111112249bbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd151:mariog=956'hfffffffffffffffffffffffffffffffffffffffe51111222129b999999999999999998888888888888872000111111111111111111111111102788889aaaaaaaaaaaaaaaaaaaa999999999aaaaabba20111111111111225abbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd152:mariog=956'hffffffffffffffffffffffffffffffffffffffffe41111222105aa999999999888888888888888888840010111111111111111111111111003888889aaaaaaaaaaaaaaaaaaaaa9999999999aaaabc601111111111112237bbbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd153:mariog=956'hfffffffffffffffffffffffffffffffffffffffffd621123221016aa9998888888888888888888886200001111111111111111111111001268888899aaaaaaaaaaaaaaaaaaa999999999999aaabba201111111111112249bacfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd154:mariog=956'hfffffffffffffffffffffffffffffffffffffffffeca7433221100159aa9988888888888888898620001111111111111111143100001247888888999aaaaaaaaaaaaaaaaaa9999999999999aaabc501111111111112237bbaefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd155:mariog=956'hffffffffffffffffffffffffffffffffffffffffffcbbbb42211110001478999999999999876300001101111111111111113667777899888888899999aaaaaaaaaaaaaa999999999999999aaabc901111111111112226ababffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd156:mariog=956'hffffffffffffffffffffffffffffffffffffffffffcbaaa522111111100001235556654321000010011111111111111111156778888888888889999999aaaaaaaaaa999999999999999999aaabb20111111111111225abbbdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd157:mariog=956'hffffffffffffffffffffffffffffffffffffffffffdbaaa8222111111110010000000000000110100111111111111111104778888886578888999999999aaaaaaa99999999999999999999aabc501111111111112249bbacfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd158:mariog=956'hffffffffffffffffffffffffffffffffffffffffffecaaaa51211111110011111101000011011101111111111111111103778888887557888999999999a99aaaa999999999999999999999aac80111111111112236abbabffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd159:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffdbaaa9311111111001111010101001011111111111111111111113788888986567788899999999999a9a99999999999999999999999aba1011111111122347abbabfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd160:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffebbaaa8111111110011111110111111111111111111111111100588889997557788889999999999999999999999999999999999999abc3011111111222479bbbabefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd161:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffdbaaaa721111111100111111111111111111111111111110137888898755788888999999999999999999999999999999998899999ab30111111223357abbbaacfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd162:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffebbaaaa8311111100352111111111110102553210000011478888987556788899999999999999999999999999999999988888899ab4122233344579abbbaabdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd163:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffdbaaaaaa62100137986111111111111036677777666678988898755678889999999999999999999999999999999998888888889a53455544448bbbbbaabeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd164:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffcbaaaaaaa98899988873111111110158777888888888888875557889999999999999999999999999999999999988888888889944565422224abbaabceffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd165:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffebbaaaaa999999988888631000014667888888888887765556789999999999999999999999999999999999998888888888898444543322236bbbdefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd166:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffdbaaaaaa9999999888899866678877655566665555556788999999999999999999a999999999999999999888888888888873344433222249babfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd167:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffdbaaaaaaa99999999888888888888877767777788899999999999999999999999999999999999999999888888888888853333333222249bbbdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd168:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffcbaaaaaa999999999998888888888888999999aaaaaaaaaa999999999999999999999999999999998888888888878742333333323348bbacffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd169:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffcbaaaaa999999999999999999999999aaaaaaaaaaaaaa9999999999999999999999999999999998888888888778721222222223347bbbbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd170:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffcbaaaaa99999999999999999999999aaaaaaaaaaaa999998888899999999999999999999999888888888877785111111223333333369efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd171:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffcbaaa999999999999999999999999aaaaaaaaa999998888888999999999999999999999999888888887777730111222333333333323bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd172:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffcbaaa999999999999999999999999999999999988888888999999999999999999999999888888887777762011112333332111122322bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd173:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffcbaaa999999999999999999999999999998888888888999999999999999999999999988888887777774111112233321000000002335cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd174:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffdbaa9999999999999999999999998888888888888999aa99aa999999999999999988888888777777301111223332000000000000124affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd175:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffcaaa99999999999999999999999988888899999aaaaaa9aa999999999999999888888887777751011212333200000000000000000137cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd176:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffebaa999999999999999999999999999999a9aaaaaaaa9a9999999999999988888887777776201112123332000000000000000000001259effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd177:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcaaa9999999999999999999999999aaaaaaaaaaaaa9a999999999999988888887777774111112223331000000000000000000000011248effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd178:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcaaa99999999999999999999999aaaaaaaaaaa9a9999999999999888888877777762011122223331000000000000000000000000011227dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd179:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecaa9999999999999999999a99a9aaaaaaaa9a9999999999999888888877777731111122223331000000000000000000000000000111235cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd180:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecba99999999999999999aaaaaaaaaa9a999999999999999888888777777520111222223331000000000000000000000000000001111226cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd181:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa54699999999999999999999999999999999999999998888887777776311112222223331000000000000000000000000000000000111226dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd182:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd744434799999999999999999999999999999999999988888887777764111122222223332000000000000000000000000000000000000111237effffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd183:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa54444441289999999999999999999999999999999988888887777775211122222222333200000000000000000000000000000000000000011124afffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd184:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd744443440000389999999999999999999999999988888888777777752112222222222333300000000000000000000000000000000000000000011124bfffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd185:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeb8544444531110012699999999999999999999988888888887777666531112222222222333310000000000000000000000000000000000000000000011227dfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd186:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffd85554444452111002210289888898998989898888888888877777666631112222222222223332000000000000000000000000000000000000000000000011123bffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd187:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffb633665554441111002211000488888888888888888888777777666665211122222222222323332000000000000000000000000000000000000000000000000011126dffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd188:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffe9533367555454211101121100000158878788888777777777766666654211122222222222232333310000000000000000000000000000000000000000000000000011124afffffffffffffffffffffffffffffffffffffffffffffffff;
10'd189:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffc84333267665565222100121100000000257777777777776666666665421112222222222222332333320000000000000000010000000100000000000000000000000000011127ffffffffffffffffffffffffffffffffffffffffffffffff;
10'd190:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffea53322216866666532210111110000000000003566666666666655543211112222222222222323333332000000000001001000000010000000000000000000000000000000001124cffffffffffffffffffffffffffffffffffffffffffffff;
10'd191:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffe9533222225877767533310111110000000000000000123444443321000111222222222222223333333332100000000001111100000000001000000000000000000000000000000111239fffffffffffffffffffffffffffffffffffffffffffff;
10'd192:mariog=956'hffffffffffffffffffffffffffffffffffffffffffff8422221111487777763342001111000000000000000000000000000000022222222222222223333333333310000000000011100000000100100000000000000000000000000000000011126efffffffffffffffffffffffffffffffffffffffffff;
10'd193:mariog=956'hfffffffffffffffffffffffffffffffffffffffffe8322211111048777776444201111100000000000000000000000000000012222222222222233333333333332000000000001111110000000000101010000000000000000000000000000001114bffffffffffffffffffffffffffffffffffffffffff;
10'd194:mariog=956'hfffffffffffffffffffffffffffffffffffffffe94221111111028777786434201111110000000000000000000000000000012222222222233333333333334433100000000001011100000000000000010101000000000000000000000000000011239fffffffffffffffffffffffffffffffffffffffff;
10'd195:mariog=956'hffffffffffffffffffffffffffffffffffffffa4222111110002887778643420011111000000000000000000000000000000222222223233333333333344444320000000000000101100000000001010010101000000000000000000000000000011127efffffffffffffffffffffffffffffffffffffff;
10'd196:mariog=956'hffffffffffffffffffffffffffffffffffffb5222111110010178777864342001111100000000000000000000000000000023333333333333333333444444432000000000000011100000000000000010101101010000100000000000000000000001124cffffffffffffffffffffffffffffffffffffff;
10'd197:mariog=956'hffffffffffffffffffffffffffffffffffd6322111110000006877786434200111110000000000000000000000000000002333333333333333334444444454310000000000000011100000000000001010110101000000000000000000000000000001123bfffffffffffffffffffffffffffffffffffff;
10'd198:mariog=956'hffffffffffffffffffffffffffffffffe83221111000000005877787434300111111000000000000000000000000000001444444444444444444444554555320000000000000010100000000000000000101011010100100000000000000000000000001238ffffffffffffffffffffffffffffffffffff;
10'd199:mariog=956'hfffffffffffffffffffffffffffffff93211111100000000487778643430011111111000000000000000000000000012455555555555555555555555555543100000000000000000100000000000010100101111010110100000000000000000000000011127fffffffffffffffffffffffffffffffffff;
10'd200:mariog=956'hfffffffffffffffffffffffffffffb5221111100011000028888864443000111111100000000111111000000012456666656655555555555555555555555320000000000000000100000000000000000000101111010100000000000000000000000000001126efffffffffffffffffffffffffffffffff;
10'd201:mariog=956'hfffffffffffffffffffffffffffe72211111010010100018888874432000011111101010111100000001234566766666665579cddddb96556665665556653100000000000000000000000000000000010111101111010101001000000000000000000000001124dffffffffffffffffffffffffffffffff;
10'd202:mariog=956'hffffffffffffffffffffffffff9321111110000000000068888744346652111000000000001123445667766666666666648dffffffffeec955666665565420000000000000000000000000000000000000000101011011111101000100000000000000000011113cfffffffffffffffffffffffffffffff;
10'd203:mariog=956'hffffffffffffffffffffffffc622111110000000035525888874443667776655444444455666777776666666666666665bffffffffeeeeeeb75666556653100000000000000000000000000000000000000111101011110101010000000000000000000000011113bffffffffffffffffffffffffffffff;
10'd204:mariog=956'hfffffffffffffffffffffff9311111100000003aeffffc98885443566776777777777777766666666666666666666667dfffffffffeeeeeeed85665666420000000000000000000000000000000000000000001111111011101101010000000000000000000001123bfffffffffffffffffffffffffffff;
10'd205:mariog=956'hfffffffffffffffffffffc521111000000002bfffffeed8785443566776666666666666666666666666666666666667efffffffffffeeeeeeed85556653200000000000000000000000000000000000000100101111111111111101010100000000000000000001113affffffffffffffffffffffffffff;
10'd206:mariog=956'hffffffffffffffffffffb321110100000005effffffeec676443466677666666666666666666666666666666666666cffffffffffeeeeeeeeedc65566531000000000000000000000000000000000000000000001111011110111111010100000000000000000011113bfffffffffffffffffffffffffff;
10'd207:mariog=956'hfffffffffffffffffff9211111000000007fffffffeed9664434666666666666666666666666666766666666666669ffffffffffefeeeeeeeddda56664200000000000000000000000000000000000000000001001111011111111111011000000000000000000011224cffffffffffffffffffffffffff;
10'd208:mariog=956'hfffffffffffffffffe5211101000000008ffffffffeeb664443667777666666667776777766666666666666666666dffffffffffeeeeeeeeedddc756532000000000000000000000000000000000000000000000101011011111111111110000000000000000000001124dfffffffffffffffffffffffff;
10'd209:mariog=956'hffffffffffffffffe5211100000000007ffffffffeed7554435667666666666666666666666666666666666666668effffffffffeeeeeeeeedddc9565310000000000000000000000000000000000000000000000000111111111111111111101000000000000000011227effffffffffffffffffffffff;
10'd210:mariog=956'hfffffffffffffffe4210000000000004fffffffffeda554434667766666666666666666666666666666666666665affffffffffeeeeeeeeeddddca5552000000000000000000000000000000000000000000000001000001011111111111110100000000000000000111138ffffffffffffffffffffffff;
10'd211:mariog=956'hffffffffffffffd4211000000000002dffffffffeeb6544346667666666666666666666666666666666666666666bfffffffffeeeeeeeeeedddcca4542100000000000000000000000000000000000000000000000000100101101110101111001000000000000000001124bfffffffffffffffffffffff;
10'd212:mariog=956'hfffffffffffffe5211000000000000affffffffeec76544466677666666666666666667766666666666666666665afefffffffeeeeeeeeeddddcca45422000000000000000000000000000000000000000000000000000100100100000000000000000000000000000011226dffffffffffffffffffffff;
10'd213:mariog=956'hfffffffffffff71000000000000004ffffffeeeed8654446667766666666666666666666666666666666666666659eeeeeeeeeeeeeeeeeddddccba443231000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011139efffffffffffffffffffff;
10'd214:mariog=956'hffffffffffff82000000000000000bfffeeeeeed95644456676666666666666666666666666666666666666666648eeeeeeeeeeeeeeeedddddccb9333243000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011126bfffffffffffffffffffff;
10'd215:mariog=956'hfffffffffffa21000000000000003efeeeeeeeda66444566666666667666666666667766666666666666666666657deeeeeeeeeeeeeedddddccba83332450000000000000000000000000000000000000000000000000000000000000110000000000000000000000000001149effffffffffffffffffff;
10'd216:mariog=956'hffffffffffd410000000000000007feeeeeeedb6654446677666666666666666666666667666666666666666765559eeeeeeeeeeeeddddddccba962323452000000000000000000000000000000000000000000000000000000000001111000000000000000000000000001126cffffffffffffffffffff;
10'd217:mariog=956'hffffffffff610000000000000000bfeeeeeedb66644466666666666666666666666666666666666666666666666556cddeeeeeedddddddcccbb9833333555100000000000000000000000000000000000000000000000000000000011110000000000000000000000000000124aefffffffffffffffffff;
10'd218:mariog=956'hfffffffffa200000100000000002deeeeeddc7665445666666666666666666666666666666666666666666656666558dddddddddddddcccbba995233335553000000000000000000000000000000000000000000000000000000001111110000000000000000000000000001128cfffffffffffffffffff;
10'd219:mariog=956'hffffffffe4100111110000000003eeeedddc766544566666666666666666666676666776666666666666665346666558cddddddddcccccbba9962243245555100000000000000000000000000000000000000000000000000000001111110000000000000000000000000000125aeffffffffffffffffff;
10'd220:mariog=956'hffffffff91000111111000000004eeddddc76764446666666666666666666666666666666666666666666664245666557bccccccccccbbaa996224522455554000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001149cffffffffffffffffff;
10'd221:mariog=956'hfffffffe41001111111000000004dddddb85764445666666666666666666666666666666666666666666666652356666568bbccbbbbbaa99852246423455555300000000000000000000000000000000000000000000000000011111111100000000000000000000000000000128bffffffffffffffffff;
10'd222:mariog=956'hfffffff910001111111100000002cdccb7576443466666666666666666666666666666666666666666666666663246666555789aaa999985223566323555555520000000000000000000000000000000000000000000000001111111111110000000000000000000000000000127bdfffffffffffffffff;
10'd223:mariog=956'hffffffe510001111111110000000adca75654323666666666666666666666666666676666666666666666666666423566655555566654322356665323555555552000000000000000000000000000000000000000000000001111111111100000000000000000000000000000025acfffffffffffffffff;
10'd224:mariog=956'hffffffc3100011111111110000006ca756533246666666666666666666666666666666666666666666666666666652356666555544444456666665224555555555100000000000000000000000000000000000000000000111111111111110000000000000000000000000000114abfffffffffffffffff;
10'd225:mariog=956'hffffff82100011111111111000000755753225666666666666666666666666666666666666666666666666666666663246666666666666666655542345555555555100000000000000000000000000000000000000000011111111111111100000000000000000000000000000149beffffffffffffffff;
10'd226:mariog=956'hffffff51000001111111111100003777532256666666666666666666666666666666666666666666666666666666666423566666555544433333332345555555555510000000000000000000000000000000000000000111111111111111010000000000000000000000000001139beffffffffffffffff;
10'd227:mariog=956'hfffffe4100000111111111111002788532266777666666666666666666666667666666766666666666666666666666665234443333322222222222335555555555555100000000000000000000000000000000000000111111111111111110000000000000000000000000000114abdffffffffffffffff;
10'd228:mariog=956'hfffffc2100001111111111111103785323667766666666666666666666666676666676666666666666666666666666666632222222222222222222335555555555555520000000000000000000000000000000000000111111111111111110000000000000000000000000000024aadffffffffffffffff;
10'd229:mariog=956'hfffffb1100000111111111111102753236667666666666666666666666666666666666666666666666666666666666666664222223334445555555555555555555555553000000000000000000000000000000000011111111111111111100000000000000000000000000000115aadffffffffffffffff;
10'd230:mariog=956'hfffff91100000111111111111102643367766666666666666666666666666666666666666666666666666666666666666666545556666666665655655555555555555555400000000000000000000000011000000011111111111111110000000000000000000000000000000126badffffffffffffffff;
10'd231:mariog=956'hfffff81000000011111111111111222677776666666666666666666666676666666666666666666666666666666666666666666666666656656555555555555555555555552000000000000000000011110000001111111111111111100000000000000000000000000000001127baeffffffffffffffff;
10'd232:mariog=956'hfffff71100000011111111111111245777666666666666666666666666666666666666666666766666666666666666666666666666666665665555555555555555555555555410000000000000002332100000011111111111111111000000000000000000000000000000001239bbeffffffffffffffff;
10'd233:mariog=956'hfffff7100000001111111111111147777766666666666666666666666666666666666666666666666666666666666666666666666665665656655555555555555555455555555410000000000013443200000001111111111111111000000000000000000000000000000000115abbfffffffffffffffff;
10'd234:mariog=956'hfffff7100000000111111111111278777666666666666666666666666666666666666666666666666666666666666666666666666666666565565555555555555555545555554455311000022454332000000111111111111111110000000000000000000000000000000000127bbcfffffffffffffffff;
10'd235:mariog=956'hfffff7100000000111111111111577777666666666666666666666666666666666666666666666666666666666666666666666666666565565655555555555555555554555544444444444444442631000000111111111111111100000000000000000000000000000000001239badfffffffffffffffff;
10'd236:mariog=956'hfffff710000000011111111111178777666666666666666666666666666666666666666666666666666666666666666666666666566665655656555555555555555555544554444444444333333362000000111111111111110100000000000000000000000000000000000125bbbefffffffffffffffff;
10'd237:mariog=956'hfffff711000000001111111111487776766666666666666666666666666666666666666666666666666666666666666666666666656656556565555555555555555555555445444444444433353350000001111111111111110000000000000000000000000000000000001139bacffffffffffffffffff;
10'd238:mariog=956'hfffff81100000000111111111168776666666666666666666666666666666666666666666666666666666666666666666666666656656555555555555555555555555545454444444444433335332000001111111111111110100000000000000000000000000000000000126abbdffffffffffffffffff;
10'd239:mariog=956'hfffffa1100000000011111111277777666666666666666666666666666666666666666666666666666666666666666666666666556565565655555555555555555555554544444444444333335320000001111111111111110000000000000000000000000000000000001139bbbfffffffffffffffffff;
10'd240:mariog=956'hfffffb210000000001111111148777666666666666666666666666666666666666666666666666666666666666666666666656656666655655555555555555555555454444444444443333333530000001111111111111110000000000000000000000000000000000000126bbadfffffffffffffffffff;
10'd241:mariog=956'hfffffd210000000000111111168777666666666666666666666666666666666666666666666666666666666666666656666566565665556555555555555555555555554445444444444333223510000011111111111111100000000000000000000000000000000000001249bbbffffffffffffffffffff;
10'd242:mariog=956'hfffffe41000000000011111127877666666666666666666666666666666666666666666666666666666666666666666666666665655655555555555555555555554545445444444444324688880000011111111111111100000000000000000000000000000000000001137bbadffffffffffffffffffff;
10'd243:mariog=956'hffffff510000000000011110387776666666666666666666666666666666666666666666666666666666666666666666656656566565555555555555555555555555554544444444436ceeeee7000011111111111111111000000000000000000000000000000000001125abacfffffffffffffffffffff;
10'd244:mariog=956'hffffff72100000000001111058776666666666666666666666666666666666666666666666666666666666666666666666656566565655555555555555555555555554544444444439eedddda0000111111111111111100000000000000000000000000000000000001239bbbefffffffffffffffffffff;
10'd245:mariog=956'hffffff9210000000000111116877666666666666666666666666666666666666666666666666666666666666666666656656566565555655555555555555555555554544444444439eeeeedd4000011111111111111100000000000000000000000000000000000001128bbadffffffffffffffffffffff;
10'd246:mariog=956'hffffffc31000000000001111787666666666666666666666666666666666666666666666666666666666666666666656656566565655555555555555555555555554544444444437eeeeeeda100011111111111111110000000000000000000000000000000000001126bbabfffffffffffffffffffffff;
10'd247:mariog=956'hffffffe5110000000001110387776666666666666666666666666666666666666666666666666666666666666665666666666565565555555555555555555554554544444444435deffeeee900001111111111111110000000000000000000000000000000000001124abbbefffffffffffffffffffffff;
10'd248:mariog=956'hfffffff8110000000000010487766666666666666666666666666666666666666666666666666666666666666656666566565655555555555555555555555555545444444444439effffeee800011111111111111111000000000000000000000000000000000001239bbadffffffffffffffffffffffff;
10'd249:mariog=956'hfffffffb21100000000000058777666666666666666666666666666666666666666666666666666666666666666666566565655655555555555555555555555545454444444434cffffffffb1011111111111111110000000000000000000000000000000000001238bbacfffffffffffffffffffffffff;
10'd250:mariog=956'hfffffffe41100000000001897766666666666666666666666666666666666666666666666666666666666666566665665656556555555555555555555555555554544444444335effffffffd301111111111111111100000000000000000000000000000000001137bbabffffffffffffffffffffffffff;
10'd251:mariog=956'hffffffff7210000000005ff87766666666666666666666666666666666666666666666666666666666666666665656656565565655555555555555555555555545444444444337ffffffffffa0011111111111111100000000000000000000000000000000001127bbabeffffffffffffffffffffffffff;
10'd252:mariog=956'hffffffffc2110000002bffd87766666666666666666666566666666666666666666666666666666566666666666566565655655555555555555555555555555454444444443437fffffffffff601111111111111100000000000000000000000000000000001126bbbbefffffffffffffffffffffffffff;
10'd253:mariog=956'hffffffffe411000004efffd77666666666666666666666666666666566666666666666656666666666656566565665655556555555555555555555555555554545444444444337fffffffffffe3011111111111100000000000000000000000000000000001125abbadffffffffffffffffffffffffffff;
10'd254:mariog=956'hfffffffff82100007fffffb77666666666666656666666665656665666666565656666566665666566565665666556565565555555555555555555555555555444444444443336efffffffffffe30111111111111000000000000000000000000000000001125abbadfffffffffffffffffffffffffffff;
10'd255:mariog=956'hfffffffffc31000affffffa77666666666666656566666666566656666566656666565666656666665656656566565655656555555555555555555555555554544444444433323dffffffffffffe301111111111100000000000000000000000000000001225abbacffffffffffffffffffffffffffffff;
10'd256:mariog=956'hffffffffff6101bffffffea77666666666556666656666655556566555656666565656656566666656666565665656556555555555555555555555555555545454444333233333bfffffffffffffe4011111111100000000000000000000000000000001225abbacfffffffffffffffffffffffffffffff;
10'd257:mariog=956'hffffffffffa11bffffffee9776666665665655666556566666655656565666656566666656656565666656566565655656556555555555555555555555544433333334445444437effffffffffffff60111111100000000000000000000000000000001225abbacffffffffffffffffffffffffffffffff;
10'd258:mariog=956'hffffffffffd4cfffffeeed876666666665656656655565555555555566665656555665656666565656656566565655656555555555555555555544444343444555555544444433adeffffffffffffff801111100000000000000000000000000000001225abbacfffffffffffffffffffffffffffffffff;
10'd259:mariog=956'hfffffffffffdfffffeeedc877666666666556555555555565555555655556565556556556565656666565665656556565555655555554444434444555555555555444444434335ecdeffffffffffffffa101110100000000000000000000000000011225abbacffffffffffffffffffffffffffffffffff;
10'd260:mariog=956'hfffffffffffffffeeeedda66766666666655656655565555555565555655565565556555565656556565665656656555554444444444455556565555555555544444444434333aedbdeffffffffffffffe3010100000000000000000000000000011225abbacfffffffffffffffffffffffffffffffffff;
10'd261:mariog=956'hffffffffffffffeeeddcba75556666666565655655655555555665555565555555555655656666565655555454444444445555666666665555555555555544444444444443435deeccdeeffffffffffffff70000000000000000000000000000011225abbacffffffffffffffffffffffffffffffffffff;
10'd262:mariog=956'hffffffffffffeeeeddcba997654445555566666565655656665656565656656565655555555444444334444555656666666666665555555555555555555454444444444434338eeefccdeeffffffffffffffb10000000000000000000000000011225abbacfffffffffffffffffffffffffffffffffffff;
10'd263:mariog=956'hfffffffffffeeeedccba998777766554444444444444444444444444444444443434434444455556667676666666666665555555555555555555555545454444444444434334cefeeebbdeeeefffffffffffff700000000000000000000000001226abbacffffffffffffffffffffffffffffffffffffff;
10'd264:mariog=956'hfffffffffeeeeedcbaa9db7766666666666666555555555555555555556565666666666666666666666666666565555555555555555555555555555554545444444444443327eeefeeebbdeeeefffffffffffffc300000000000000000000001226abbacfffffffffffffffffffffffffffffffffffffff;
10'd265:mariog=956'hfffffffffeeeddcbaa9cfa766666666666666666666666666666666666666666666666666666666666556556565555555555555555555555555555554545444444444443333aeefefeeebbdeeeeeeffffffffffff9100000000000000000001125abbacffffffffffffffffffffffffffffffffffffffff;
10'd266:mariog=956'hffffffffeeeddcbaa9cffa776666666666656665566655656666656565655656565655556565655556555555555555555555555555555555555555545444544444444433334deeefeffeebacdeeeeeeeeffffffffff9100000000000000001126bbbacfffffffffffffffffffffffffffffffffffffffff;
10'd267:mariog=956'hffffffffeeddcbaaabfffa766666565556555555556555555556555655555555555555555555555555555555555555555555555555555555555555454544444444443333326eeefeffffeebacddeeeeeeeeeefffffffe9200000000000000124abbacffffffffffffffffffffffffffffffffffffffffff;
10'd268:mariog=956'hffffffffeddcbaaaaffffa766666565555555555565555555555555555555555555555555555555555555555555555555555555555555555554554444444444333333333329eeeffffffffebabcddeeeeeeeeeeefffffffa4000000000001138abbdfffffffffffffffffffffffffffffffffffffffffff;
10'd269:mariog=956'hffffffffedcbaaaaeffffa77666666655555555555555555555555555555555555555555555555555555555555555555555555555555545454444444443433344445543333ceefffffffffffcabcddddeeeeeeeeeeeeffffffa4000000000379abbefffffffffffffffffffffffffffffffffffffffffff;
10'd270:mariog=956'hfffffffffdcbaaaefffff966666665555555555555555555555555555555555555555555555555555555555555555555555555545444444444344444445555555444543335deeffffffffffffdaabcdddddddedeeeeeeeeeefffeb8431125899abbbfffffffffffffffffffffffffffffffffffffffffff;
10'd271:mariog=956'hfffffffffdbaaacffffff956666555555555555555555555555555555555555555555555555555555555555555555555555444443343444455555555555544444444543326eeefffffffffffffdaabbcddddddddddddeeeeeeeeffffffffeedcbbcbdffffffffffffffffffffffffffffffffffffffffff;
10'd272:mariog=956'hfffffffffebaaafffffffb65555555555555555555555555555555555555555555555555555555555555555555444444444444555556655555554544444444444444534338eeefffffffffffffffbaabbcccddddddddddddeeeeeeeeeeeeeeeeedcbbffffffffffffffffffffffffffffffffffffffffff;
10'd273:mariog=956'hffffffffffcaadfffffffb8765455555555555555555555555555555555555555555555555555555444444444444545556665555555555545444544444444444444453333aeeeffffffffffffffffc9abbbccccccccccddddddeeeeeeeeeeeeeddcbbefffffffffffffffffffffffffffffffffffffffff;
10'd274:mariog=956'hfffffffffffbcffffffffc6777765444444555555555555555555555555555545444444444444444545555666666665555555554555555454545444444444444444333333beeefffffffffffffffffd99ababbcccccccccccccddddddeeeedddcccbaefffffffffffffffffffffffffffffffffffffffff;
10'd275:mariog=956'hfffffffffffffffffffffc7665666766655544444444444444444444444444444455555566666666666665555555555555555555555554445444444444444444444443334ceeffffffffffffffffffffb88aaaabbbbbbbbbbbbccccccccccccbbcbbbefffffffffffffffffffffffffffffffffffffffff;
10'd276:mariog=956'hfffffffffffffffffffffd7666555555566666666666666666666666666666666666666655555555555555555555555555555555545444544444444444444444443443335deeeffffffffffffffffffffea89aaaaaabbbbbbbbbbbbbbbbbbbbbbbbbbefffffffffffffffffffffffffffffffffffffffff;
10'd277:mariog=956'hfffffffffffffffffffffe7666555555555555555555566555555555555555555555555555555555555555555555555555555555454445444444444444444444443433326deeeffffffffffffffffffffffc989aaaaaaaaaaaaaaababbbbbbbbbbbbbffffffffffffffffffffffffffffffffffffffffff;
10'd278:mariog=956'hffffffffffffffffffffff8666665555555555555555565555555556555555555555555555555555555555555555555555555554544444444444444444444444433433327deeefffffffffffffffffffffffea8889aaaaaaaaaaaaaaaaaaabbbbbbacffffffffffffffffffffffffffffffffffffffffff;
10'd279:mariog=956'hffffffffffffffffffffffa666655555555555555555555555555555555555555555555555555555555555555555555555555544444444444444444444444444433443328deeeffffffffffffffffffffffeeeb987899aaaaaaaaaaaaaaaaabcbbbbeffffffffffffffffffffffffffffffffffffffffff;
10'd280:mariog=956'hffffffffffffffffffffffb666655555555555555555556555555555555555555555555555555555555555555555555555554545444444444444444444444444333443329eeeeffffffffffffffffffffffeeeec98778999aaaaaaaaaaaaabbcbbadfffffffffffffffffffffffffffffffffffffffffff;
10'd281:mariog=956'hffffffffffffffffffffffc666555555555555555555566555555555555555555555555555555555555555555555555555545444444444444444444444444443333343329deeeffffffffffffffffffffffeeeddb98888889999aaaaaaaabbbccbcffffffffffffffffffffffffffffffffffffffffffff;
10'd282:mariog=956'hffffffffffffffffffffffd76665555555555555555555555555555555555555555555555555555555555555555555545544444444444444444444444444443433334432aeeeeffffffffffffffffffffffeeeddca99998888899999aaaabbbccbcffffffffffffffffffffffffffffffffffffffffffff;
10'd283:mariog=956'hffffffffffffffffffffffe86655555555555555555555655555555555555555555555555555555555555555555555554454444444444444444444444444333333333343aeeeefffffffffffffffffffffeeeeddcbaa99999999999aaaabbbbccbbffffffffffffffffffffffffffffffffffffffffffff;
10'd284:mariog=956'hfffffffffffffffffffffffa6655555555555555555555555555555555555555555555555555555555555555555555444444444444444444444444444444433333333323beeeefffffffffffffffffffffeeeeddcbaaaa999999aaaaaaabbbbccbaefffffffffffffffffffffffffffffffffffffffffff;
10'd285:mariog=956'hfffffffffffffffffffffefb6655555555555555555555655555555555555555555555555555555555555555555454444444444444444444444444444444333333333322beeeefffffffffffffffffffffeeeeddcbaaaaaaaaaaaaaaaaabbbbbccadfffffffffffffffffffffffffffffffffffffffffff;
10'd286:mariog=956'hffffffffffffffffffffeeee7655555555555555555555555555555455555555555555555555555555555555554444444444444444444444444444443443333333333322bdeeeefffffffffffffffffffeeeeeddcbaaaaaaaaaaaaaaaaabbbbbccacfffffffffffffffffffffffffffffffffffffffffff;
10'd287:mariog=956'hfffffffffffffffffffeeeef9665555555555555555555555555554555555555555555555555555555555545444444444444444444444444444444443433333333333222beeeeeffffffffffffffffffeeeeedddcbbbaaaaaaaaaaaaaaabbbbbccbbfffffffffffffffffffffffffffffffffffffffffff;
10'd288:mariog=956'hffffffffffffffffffeeeeefb655555555555555555555555555555555555555555555555555555555555454444444444444444444444444444444444433333333333222bdeeeefffffffffffffffffeeeeeedddcbbbaaaaaaaaaaaaaaabbbbbccbbfffffffffffffffffffffffffffffffffffffffffff;
10'd289:mariog=956'hffffffffffffffffeeeeeeeed765555555555555555555555555555455455545555545555555555545445444444444444444444444444444444433333333333333322222bdeeeefffffffffffffffffeeeeeeddccbbbaaaaaaaaaaaaaaaabbbbbcbbeffffffffffffffffffffffffffffffffffffffffff;
10'd290:mariog=956'hffffffffffffffffeeeeeeeeea65555555555555555555455555545455545454555455544545545444444444444444444444444444444444444443433333333332333333adeeeefffffffffffffffeeeeeeeeddccbbbaaaaaaaaaaaaaaaaabbbbccadffffffffffffffffffffffffffffffffffffffffff;
10'd291:mariog=956'hffffffffffffffffeeeeeeeeec76555555555555555555455454454445454545444545545444444444444444444444444444444444444444433333333333333333444444adeeeeffffffffffffffeeeeeeeedddcbbbbbbaaaaaaaaaaaaaaabbbbccbcffffffffffffffffffffffffffffffffffffffffff;
10'd292:mariog=956'hfffffffffeefeeeeeeeeeeeeee96555555555554554554455444544455445454445444454444444444444444444444444444444444444434443433334333334445555554adeeeeeffffffffffffeeeeeeeeedddcbbbbbbaaaaaaaaaaaaaaabbbbbcbbffffffffffffffffffffffffffffffffffffffffff;
10'd293:mariog=956'hfffffffffeefefeeeeeeeeeeeec65555555555545545444554444444454444444444444444444444444444444444444444444444444433344333333334444455555555549deeeeefffffffffffeeeeeeeeeeddccbbbbbbbaaaaaaaaaaaaaabbbbbccbefffffffffffffffffffffffffffffffffffffffff;
10'd294:mariog=956'hfffffffffeeeeeeeeeeeeeeeeee86555555555445444455454544444454444444444444444444444444444444444444444444434433433343433433444444555555555549ddeeeefffffffffeeeeeeeeeeedddccbbbbbbbaaaaa9aaaaaaaaabbbbbcbdfffffffffffffffffffffffffffffffffffffffff;
10'd295:mariog=956'hfffffffffeeeeeeeeeeeeeeeeeeb6555455455455445444455444444454444444444444444444444444444444444444444444433433333333334334444455555555555547ddeeeeeefffffefeeeeeeeeeeedddcbbbbbbbbaaaa999999aaaaaabbbbcbcfffffffffffffffffffffffffffffffffffffffff;
10'd296:mariog=956'hffffffffffeeeeeeeeeeeeeeeeed8655554544444444444455444444455444444444444444444444444444444444444444343334334333333443444445555555555555547cdeeeeeefffffeeeeeeeeeeeedddccbbbbbbbbaaaa9999999aaaaaabbbccbfffffffffffffffffffffffffffffffffffffffff;
10'd297:mariog=956'hfffffffffeeeeeeeeeeeeeeeeeeeb655444444444444444445444444445444444444444444444444444444444444444343443333333333344344445555555555555555546cdeeeeeeefeefeeeeeeeeeeeedddccbbbbbbbbaaa99999999aaaaaaabbbcbdffffffffffffffffffffffffffffffffffffffff;
10'd298:mariog=956'hffffffffffeeeeeeeeeeeeeeeeeed755554444544444444445444444445444444444444444444444444444444444444433333333333333434444545555555555555555555bdeeeeeeeeeeeeeeeeeeeeeedddccbbbbbbbbbbaa999999999aaaaaaabbccbffffffffffffffffffffffffffffffffffffffff;
10'd299:mariog=956'hffffffffffeeeeeeeeeeeeeeeeeeeb65544444444444444445544444444444444444444444444444444444444444444333333333333333444445555555565555555555545addeeeeeeeeeeeeeeeeeeeeedddccbbbbbbbbbbaa9999999999aaaaaabbbcbefffffffffffffffffffffffffffffffffffffff;
10'd300:mariog=956'hffffffffffeeeeeeeeeeeeeeeeeedd855545444444444444445444444445444444444444444444444444444444444333333333333333444445555555556556555555555548ddeeeeeeeeeeeeeeeeeeeeeddccbbbbbbbbbbaaaa999999999999aaaabbcccfffffffffffffffffffffffffffffffffffffff;
10'd301:mariog=956'hffffffffffeeeeeeeeeeeeeeeeeedec65444444444444444445444444435444444444444444444444444444444343333333333333334444555555565565565555555555547cdeeeeeeeeeeeeeeeeeeeedddccbbbbbbbbbbaaa9999999999999aaaabbbcbdffffffffffffffffffffffffffffffffffffff;
10'd302:mariog=956'hffffffffffeeeeeeeeeeeeeeeeeeddd95544444444444444444545545444444444444444444444444444444443333333333333334444445555555655655655555555555546cdeeeeeeeeeeeeeeeeeeedddccbbbbbbbbbbaaaa99988888889999aaaabbbcbffffffffffffffffffffffffffffffffffffff;
10'd303:mariog=956'hfffffffffffeeeeeeeeeeeeeeeeedddc7554444444444444444544443444444444444444444444444444444333333333333333334444555555556555556656655555555545bddeeeeeeeeeeeeeeeeeedddcbbbbbbbbbbaaaaa999888888889999aaabbbcbdfffffffffffffffffffffffffffffffffffff;
10'd304:mariog=956'hfffffffffffeeeeeeeeeeeeeeeeeddddb6544444444444444444434344434444444444344444444444344333333333333333334444455555555655665655665555555555549ddeeeeeeeeeeeeeeeeedddccbabbbbbbbaaaaa999ba88888889999aaabbbbcbfffffffffffffffffffffffffffffffffffff;
10'd305:mariog=956'hfffffffffffeeeeeeeeeeeeeeeeeddddd9554444444434344444544434333534443444434344343433333333333333333333344444555555556556556656655555555555548ddeeeeeeeeeeeeeeeedddccbbbbbbbbbaaaaa999ab987778889999aaaabbbcccffffffffffffffffffffffffffffffffffff;
10'd306:mariog=956'hfffffffffffeeeeeeeeeeeeeeeeeddddcb754444444434433433543344433443433343333333334333333333333333333333444455555555555566566556565555555555546cdeeeeeeeeeeeeeeedddccbbabbbbaaaaaaa9999bba777778889999aaaabbbcbefffffffffffffffffffffffffffffffffff;
10'd307:mariog=956'hffffffffffffeeeeeeeeeeeeeeedddddcca65444444434333333353333333344333333333333333333333333333333333333444555555555655665665665565655555555555bddeeeeeeeeeeeeedddccbaabbbbbaaaa999999abac989987788899aaaabbbbccfffffffffffffffffffffffffffffffffff;
10'd308:mariog=956'hfffffffffffeddeeeeeeeeeeeeeddddcccb65554444433433333345333333343333333333333333333333333333333333344445555555555556655655655656655555555544addeeeeeeeeeeeedddccbaaaabbbaaaa9999999aabefffffeb889999aaaabbbbccffffffffffffffffffffffffffffffffff;
10'd309:mariog=956'hffffffffffeeddeeeeeeeeeeeeeeddddccb855554444344333333344333333343333333333333333333333333333333333444555555555555665665565565565555555555548cddeeeeeeeeeedddccbaaaaabaaaa999888999acfffffffffc89aaaaaaabbbbcbdfffffffffffffffffffffffffffffffff;
10'd310:mariog=956'hfffffffffeedccdeeeeeeeeeeeeddddcccb955444544444443433335333333334333333333333333333333333333333334455555555555556655665655655656555555555546bddeeeeeeeeedddccbaaaaabaaaa99888888989fffffffffffc99aabaaaabbbbcbfffffffffffffffffffffffffffffffff;
10'd311:mariog=956'hffffffffeeddefedeeeeeeeeeeeddddccbba65454444444444333333533333334433333333333333333333333333333344555555555566556556656656556555555555555544addeeeeeeeedddccbaaaaaaaaaaa9877777887cfffffffffeed99aabbaaaabbbcbcffffffffffffffffffffffffffffffff;
10'd312:mariog=956'hfffffffeedeffffddeeeeeeeeeeddddccbbb654444454444443343333533333334333333333333333333333333333334445555555555555665565665665655655555555555548cddeeeeeeddddccbaaaaaaaaa998776666779efffffffffedcbcdddcbaaaabbbbbefffffffffffffffffffffffffffffff;
10'd313:mariog=956'hfffffffeffffffffddeeeeeeeeddddccbbba755444444444444434333353333333533333333333333333333333333334555555555555555655656666656656555555555555545bddeeeedddddccbbababaaaa998766556677cfffffffffeedbdeeeedcaaaaabbbadfffffffffffffffffffffffffffffff;
10'd314:mariog=956'hffffffefffffffffedeeeeeeeeddddccbbaa8554444444444434334333443333333533333333333333333333333333445555555555555565566566665665665555555555555449cdddedddddccbbaaaaaaa99887655555668effffffffeedcbdfeeecba9aaaabbbbfffffffffffffffffffffffffffffff;
10'd315:mariog=956'hffffffffffffffffffeeeeeeeedddccbbaa97555444444444333333333344333333343333333333333333333333334455555555555555665665565665656656555555555555546cddddddddccbbaaaaaaa87776654445557affffffffeedcbbbdedcbba9aaaabbbbeffffffffffffffffffffffffffffff;
10'd316:mariog=956'hfffffeeffffffffffffeeeeeedddccbba99875555444344434333333333334333333433333333333333333333333445555555555555565556566566565565655555555555555449cdddddddcbaaaaaabbb96555664334567cfffffeeeedcbbb9acbaab9999aabbbbeffffffffffffffffffffffffffffff;
10'd317:mariog=956'hfffffeeeeffffffffffeeeeedddccbba988775555444333433333333333333333333333333333333333333333333444555555555555555565565565665655556555555555555545bddddddccbbbbbbbbaab9678887546668effffeeeeddcbba99aaaba899aabbbbbfffffffffffffffffffffffffffffff;
10'd318:mariog=956'hfffffedeeeeffffffffeeeeddddccba98887765555443333333333333333333333333333333333323333333334334445555555555555555656556566566565655555555555554447ddddddddddeeeeeedbaa87888767776aefffeeeeddcbaba99aaaa999aabbbbadfffffffffffffffffffffffffffffff;
10'd319:mariog=956'hffffffdddeeeeeeeeeeeeeddddcbba988877665555543433333333333333233333333333333333322222233334334555555555555555556555565565655656555555555555554544adddddeeeeeeeeeeedb977888677888bffffeeeddcbaab99aaabbbbbbbbbaacffffffffffffffffffffffffffffffff;
10'd320:mariog=956'hfffffffccddeeeeeeeeedddddcba998887776655555543333333333333322222233333323333333222222233334345455555555555555655656656566565565655555555555554446cdddeeeeeeeeeeeedddca88777888aeeffeeeedccbaba99aaabbbbaaaabcefffffffffffffffffffffffffffffffff;
10'd321:mariog=956'hfffffffebcdddddddddddcccba99988887776655555544333333333333333222212222323222223222222233334445555555555555555556556565565665656555555555555554444adddeeeeeeeeeeeefffffec76778aefeeeeedddcbaab99aaabbbabccdeffffffffffffffffffffffffffffffffffff;
10'd322:mariog=956'hffffffffebbccdddccccbbaa99999888877788655555544333333333333333222222222222222222222222333334555555555555555555555655656556565655555555555555554445bdddeeeeeeeeeeffffffffdbefffffeeeedddcbaaaa9aaaabbbbeffffffffffffffffffffffffffffffffffffffff;
10'd323:mariog=956'hfffffffffebabbcccbbaa999999988888888886555555544333333333333333322222222222222222222223333344555555555555555555556565665656556565555555555555444447cddeeeeeeeefffffffffffffffffffeedddcbbaaa9aaaaaaabdfffffffffffffffffffffffffffffffffffffffff;
10'd324:mariog=956'hffffffffffebaaaaaa9999999999999998888876555555554333333333333333332222222222222222222223333455555555555555555555556556565665656555555555555555544438cddeeeeeeeffffffffffffffffffffedcccaaaaa9aaaa99aaefffffffffffffffffffffffffffffffffffffffff;
10'd325:mariog=956'hffffffffffffcaaaa99999999aaa998888889a86655555555433333333333333332222222222222221111112333455555555555555555555556566665656565555555555555555454443acddeeeeefffffffffffffffffffffeecbaaaaa99aaa9899aadffffffffffffffffffffffffffffffffffffffff;
10'd326:mariog=956'hfffffffffffffdbaaaaaaaaaabbbaa9999aaab965555555555443333333333333332222222222222221111113334555555555555555555555656656565665655565555555555555444434acdddeeeeffffffffffffffffffffeecaaaaa999aa98999aabdfffffffffffffffffffffffffffffffffffffff;
10'd327:mariog=956'hfffffffffffffffdbabbbbbbbbaaaabbbbbbbba755555555555443333333333333333232222222222221111123345555555555555555556555565665556565655555555555555555544424bcdddeeeeffffffffffffffffffeeeda9aa9999a98999aaaaadffffffffffffffffffffffffffffffffffffff;
10'd328:mariog=956'hfffffffffffffffffecbbaabbbcdeecbaaaabbc8655555555555443333333333333332222222222222221111123455555555555555555555555566565656655555655555555555554444415bccdddeeeefffffffffffffffeeeedb9a99999888999aaaaabdfffffffffffffffffffffffffffffffffffff;
10'd329:mariog=956'hfffffffffffffffffffffeeeffffffffeeeefff95555555555555444333333333333332222222222222211111134455555555555555555555555656565565656565555555555555554444315abccddeeeeeefffffffffeeeedddcba999997888999aaaabbbdffffffffffffffffffffffffffffffffffff;
10'd330:mariog=956'hfffffffffffffffffffffffffffffffffffffffa665555555555555443333333333332322222222222222111112344555555555555555555555655556565655555555555555555555454442149bbcddddeeeeeeeeeeeeeeddddcbb999977888999aaaaabbbbefffffffffffffffffffffffffffffffffff;
10'd331:mariog=956'hfffffffffffffffffffffffffffffffffffffffa6655555555555555443333333333333222222222222222111112455555555555555555555555565656555565655555555555555555544432127abbcddddeeeeeeeeeddddccbbba9877778889999aaaabbbbbfffffffffffffffffffffffffffffffffff;
10'd332:mariog=956'hfffffffffffffffffffffffffffffffffffffffb665555555555555554433333333332332222222222222111111134455555555555555555555555555566565656555555555555555544444321159abbccddddddddddcccbbbaaa76677788888999aaaabbbbaeffffffffffffffffffffffffffffffffff;
10'd333:mariog=956'hfffffffffffffffffffffffffffffffffffffffd76555555555555555554433333333332222222222222222111112445555555555555555555555565656565655656555555555555555454442221269aabcccccccccbbbaaaaaa766777778889999aaaabbbbadffffffffffffffffffffffffffffffffff;
10'd334:mariog=956'hfffffffffffffffffffffffffffffffffffffffe7655555555555555555544333333332322222222222222111111134555555555555555555556565555565565655555555555555555554444322221269aaaabaaaaaaaaaaaa97666677778888999aaaaabbbacffffffffffffffffffffffffffffffffff;
10'd335:mariog=956'hfffffffffffffffffffffffffffffffffffffffe766555555555555555555443333333322222222222222212111111445555555555555555555555555566565656555555555555555555454443222221369999999999999aaaa99876677778889999aaaaabbacffffffffffffffffffffffffffffffffff;
10'd336:mariog=956'hffffffffffffffffffffffffffffffffffffffff8555555555555555555555544333333322222222222222221111112455555555555555555555556555656565655556555555555555555454442222222124789999999abbbbbbbba9877777788899aaaaabbacffffffffffffffffffffffffffffffffff;
10'd337:mariog=956'hffffffffffffffffffffffffffffffffffffffff966555555555555555555554443333323222222222222221111111254555555555555555555555555556656565656555555555555555554444322222222222336abbbbbbaabcdcbbaa987777888999aaabbacffffffffffffffffffffffffffffffffff;
10'd338:mariog=956'hffffffffffffffffffffffffffffffffffffffffa665555555555555555555554443333322222222222222212111112445555555555555555555555655565656565555555555555555555545444322222222222349bbaaabcdfffffedbaaa9888888999abbbadffffffffffffffffffffffffffffffffff;
10'd339:mariog=956'hffffffffffffffffffffffffffffffffffffffffb555555555555555555555555444333322222222222222221211112434555555555555555555555555556566555656555555555555555554444432223222333348aceeffffffffffffedbabaaaaaaabbbbabfffffffffffffffffffffffffffffffffff;
10'd340:mariog=956'hffffffffffffffffffffffffffffffffffffffffc666555555555555555555555444443323222222222222222111112324555555555555555555555555566565556565555555555555555555544442222322333346acfffffffffffffffffecbbabbbbbbaacffffffffffffffffffffffffffffffffffff;
10'd341:mariog=956'hffffffffffffffffffffffffffffffffffffffffd6655555555555555555555545444443322222222222222221212214235555555555555555555555555655565655555555555555555555554544432333333333459bffffffffffffffffffffedcbbbbbcefffffffffffffffffffffffffffffffffffff;
10'd342:mariog=956'hffffffffffffffffffffffffffffffffffffffffe7665555555555555555555554544444332222222222222222221113224555555555555555555555555566666656565555555555555555555454543322333333348bdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd343:mariog=956'hffffffffffffffffffffffffffffffffffffffffe7655555555555555555555545454444433222222222222222222213213555555555555555555555555555656565655555555555555555555555444333333333346acffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd344:mariog=956'hfffffffffffffffffffffffffffffffffffffffff7665555555555555555555554544444443322222222222222221213312455555555555555555555565656565556656555555555555555555555454433333333445abffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd345:mariog=956'hfffffffffffffffffffffffffffffffffffffffff86655555555555555555555554544444443322222222222222121133123555555555555555555555555665555565656565555555555555555555444333333334459befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd346:mariog=956'hfffffffffffffffffffffffffffffffffffffffff96655555555555555555555554544444443332222222222222222133122455555555555555555555555555565656565555555555555555555555454433333333457acfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd347:mariog=956'hfffffffffffffffffffffffffffffffffffffffffa6555555555555555555555545544444444333222222222222222134122455555555555555555555555565666565565556555555555555555555545443333333346abfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd348:mariog=956'hfffffffffffffffffffffffffffffffffffffffffb66555555555555555555555544444444444333222222222222222231222455555555555555555555556555556656565655555555555555555555555443333334459beffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd349:mariog=956'hfffffffffffffffffffffffffffffffffffffffffc66555555555555555555555554544444444433322222222222222231222455555555555555555555556565556565655555555555555555555555555444333334458adffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd350:mariog=956'hfffffffffffffffffffffffffffffffffffffffffd66555555555555555555555545444444444443332222222222222242222345555555555555555555555555565656655565655555555555555555554545433334446acffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd351:mariog=956'hfffffffffffffffffffffffffffffffffffffffffe765555555555555555555555545444444444443332222222222222322223455555555555555555555555555556555655565555555555555555555555444433344459befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd352:mariog=956'hfffffffffffffffffffffffffffffffffffffffffe756555555555555555555555554444444444444333222222222222322222355555555555555555555555656565556565655555555555555555555554544433344458bdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd353:mariog=956'hffffffffffffffffffffffffffffffffffffffffff856555555555555555555555554444444444444333222222222222422222345555555555555555555555555656565565556565555555555555555555554543334457bcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd354:mariog=956'hffffffffffffffffffffffffffffffffffffffffff9555555555555555555555555454444444444444333222222222223222222355555555555555555555555565665656565656555555555555555555555454444344459bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd355:mariog=956'hffffffffffffffffffffffffffffffffffffffffff9665555555555555555555555554444444444444433322222222224222222345555555555555555555555655656565656556555655555555555555555554444344458beffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd356:mariog=956'hffffffffffffffffffffffffffffffffffffffffffa656555555555555555555555554544444444444433332222222223222323345555555555555555555555555565656556565655555555555555555555544444444457acffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd357:mariog=956'hffffffffffffffffffffffffffffffffffffffffffb6655555555555555555555555454444444444443333332222222232222223345555555555555555555555556665565656565555555555555555555555555454434469bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd358:mariog=956'hffffffffffffffffffffffffffffffffffffffffffc6655555555555555555555545544444444444434333332222222243222223345555555555555555555555556565656565555655555555555555555555554444444458befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd359:mariog=956'hffffffffffffffffffffffffffffffffffffffffffc6555555555555555555555555544444444444444433333222222233222232345555555555555555555555565656555665556555555555555555555555554444444447adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd360:mariog=956'hffffffffffffffffffffffffffffffffffffffffffd75655555555555555555555554544444444444443333333222222332223233345555555555555555555556556655666565656555555555555555555555554544444459cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd361:mariog=956'hffffffffffffffffffffffffffffffffffffffffffe75655555555555555555555555454444444444443333333322222332222223345555555555555555555555565656565656555555555555555555555555555444444458beffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd362:mariog=956'hffffffffffffffffffffffffffffffffffffffffffe76655555555555555555555555444444444444444333333322222332222333344555555555555555555555656566656566565556555555555555555555555544455556adffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd363:mariog=956'hfffffffffffffffffffffffffffffffffffffffffff855555555555555555555555545444444444444443433333322223322222333445555555555555555555555656655565656565655555555555555555555545454555459cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd364:mariog=956'hfffffffffffffffffffffffffffffffffffffffffff966555555555555555555555554544444444444444333333332223322222233445555555555555555555555555565656565555655555555555555555555555545555547befffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd365:mariog=956'hfffffffffffffffffffffffffffffffffffffffffff965555555555555555555555555444444444444443333333333222322222333454555555555555555555656565656565565656565655555555555555555555544454556acfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd366:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffa555555555555555555555555554444444444444443333333332223222223334555555555555555555555556666556656565656555565555555555555555554545554559bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd367:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffb665555555555555555555555545544444444444443333333333223222222334564555555555555555555655655556565666655555555555555555555555555554555557aeffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd368:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffb5655555555555555555555555545444444444444443333333332232222333345855555555555555555555656565656566565556565555555555555555555555545555569cffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd369:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffc6555555555555555555555555554444444444444443333333333242222233345864555555555555555555565656566665656565555555555555555555555555554555558befffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd370:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffc6655555555555555555555555555444444444444433333333333232222232345884555555555555555555555555565656565665656555555555555555555555454555557adfffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd371:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffd66555555555555555555555555554444444444443433333333332432222333458a55555555555555555555665656566656555565655555555555555555555555555555559cfffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd372:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffd66555555555555555555555555545444444444444333333333332432222233347b65555555555555555555556565656666565656556555555555555555555555555555558beffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd373:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffe76555555555555555555555555454444444444444433333333332332222233357b85555555555555555555566665556565655555565555555555555555555555555555557acffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd374:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffe76555555555555555555555555554444444444444333333333333532222233347b955555555555555555555555555656565665656555555555555555555555555555555569bffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd375:mariog=956'hffffffffffffffffffffffffffffffffffffffffffff76655555555555555555555555554444444444444433333333333443222333346bb74555555555555555555565656566565656565565555555555555555555555555555557aefffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd376:mariog=956'hffffffffffffffffffffffffffffffffffffffffffff86655555555555555555555555554544444444444433333333333442332333346ab945555555555555555556566555656566555655655555555555555555555555555555569cfffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd377:mariog=956'hffffffffffffffffffffffffffffffffffffffffffff86655555555555555555555555554444444444444433333333332443332233346abb45555555555555555555555656565665656656555555555555555555555555554555558beffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd378:mariog=956'hffffffffffffffffffffffffffffffffffffffffffff96655555555555555555555555554444444444444333333333333443332233345abc55555555555555555555655565565656656566565555555555555555555555555555557adffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd379:mariog=956'hffffffffffffffffffffffffffffffffffffffffffff96655555555555555555555555554544444444443443333333333333332233345abd745555555555555555555555656566565655655555555555555555555555555555555569cffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd380:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffa66555555555555555555555555554444444444444333333333333433332333459bda45555555555555555555556566565656656556565555555555555555555555555555558aefffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd381:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffa66555555555555555555555555555444444444443333333333333433333333449bdc555555555555555555555555656566565665656656555555555555555555555555555569cfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd382:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffa66555555555555555555555555554444444444443433333333333433322333359bce655555555555555555555656556565655656656556555555555555555555555555555558bfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd383:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffb66555555555555555555555555554444444444444333333333333332233233448bcf845555555555555555555556565656656656565565555555555555555555555555555557adffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd384:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffb66555555555555555555555555554444444444444433333333333433332233348bcfa455555555555555555565655556565566665656655556555555555555555555555555569cffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd385:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffb66655555555555555555555555545444444444444433333333333433322333348bbfc555555555555555555555555565665656656656556555555555555555555555555555567befffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd386:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffc66555555555555555555555555554444444444444433333333333433322233447abfe645555555555555555555555555655656656556556555555555555555555555555555566acfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd387:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffc66555555555555555555555555454444444444444433333333334433322333347abff8455555555555555555555556566565665665665655555555555555555555555555555569bfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd388:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffc65655555555555555555555555554444444444444443333333333433322233447abefb455555555555555555555555565665656656655656656555555555555555555555555568adffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd389:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffc76555555555555555555555555544444444444444433333333333333233323346abefd4555555555555555555555556556566566566566565555555555555555555555555555579cffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd390:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffb666555555555555555555555555544444444444444433333333334333232333469beff6455555555555555555555556565566665565665665555555555555555555555555555568befffffffffffffffffffffffffffffffffffffffffffffffff;
10'd391:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffb665555555555555555555555555444444444444444434333333333332323323469bdff8455555555555555555555555565666655665665655655655555555555555555555555567adfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd392:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffa666655555555555555555555555554444444444444343333333344322223333459bdffb4555555555555555555555556556566566666566556565565555555555555555555555569bfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd393:mariog=956'hffffffffffffffffffffffffffffffffffffffffffff9666655555555555555555555555544444444444444433333333333333323333458bcffe5455555555555555555555555566566566566665566565565555555555555555555555568beffffffffffffffffffffffffffffffffffffffffffffffff;
10'd394:mariog=956'hffffffffffffffffffffffffffffffffffffffffffff8666666556555555555555555555544444444444444433333333344233233233458bcfff8455555555555555555555565565665666665666566566565555555555555555555555557acffffffffffffffffffffffffffffffffffffffffffffffff;
10'd395:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffd7666666666666555565555555555554444444444444443333333333332333233457abfffb4555555555555555555555556656666656656666656655655555555555555555555555569befffffffffffffffffffffffffffffffffffffffffffffff;
10'd396:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffc6666666666666665655555555555544444444444444433333333344333232233347abfffd5455555555555555555555555556556566566656656656655655555555555555555555568adfffffffffffffffffffffffffffffffffffffffffffffff;
10'd397:mariog=956'hfffffffffffffffffffffffffffffffffffffffffff97776666666666656655555555555544444444444444443333333343332333233446abefff74555555555555555555555555655656666665666566566566555555555555555555555569bfffffffffffffffffffffffffffffffffffffffffffffff;
10'd398:mariog=956'hffffffffffffffffffffffffffffffffffffffffffc76666666666666666655555555555554444444444444444333333343333333333456abefffa4555555555555555555555555656656666655665665665566555555555555555555555567aeffffffffffffffffffffffffffffffffffffffffffffff;
10'd399:mariog=956'hfffffffffffffffffffffffffffffffffffffffffd8766666666666666666555555555555544544444444444443433333433333333333569bdfffd44555555555555555555565565566566566566656656655665555555555555555555555569cffffffffffffffffffffffffffffffffffffffffffffff;
10'd400:mariog=956'hffffffffffffffffffffffffffffffffffffffffc76666666666665566666655555555555555444444444444434333333433333333333459bdffff64555555555555555555555555665665666566556656655665565555555555555555555568befffffffffffffffffffffffffffffffffffffffffffff;
10'd401:mariog=956'hfffffffffffffffffffffffffffffffffffffffc766666666666666655566665555555555545444444444444443433333433333333333458bcffff94455555555555555555655655655655665665566656655665555555555555555555555667adfffffffffffffffffffffffffffffffffffffffffffff;
10'd402:mariog=956'hffffffffffffffffffffffffffffffffffffffe7666666666666666666555665555555555554444444444444434333333433333333333457bcffffd54555555555555555555555555566556656656666666566656655555555555555555555669bfffffffffffffffffffffffffffffffffffffffffffff;
10'd403:mariog=956'hffffffffffffffffffffffffffffffffffffff96666666666666666666655565555555555555454444444444443333334433333333334456abfffff74555555555555555555555565565566566656665666566556655565555555555555555557aeffffffffffffffffffffffffffffffffffffffffffff;
10'd404:mariog=956'hfffffffffffffffffffffffffffffffffffffd66656655666666666666556555555555555545444444444444443333333433333333333446abeffffa44555555555555555555555556556656665666566655665565556655555555555555555569cffffffffffffffffffffffffffffffffffffffffffff;
10'd405:mariog=956'hfffffffffffffffffffffffffffffeeeeeeffb566555555665566666666555555555555555555444444444444443333354333333333334459beffffc54555555555555555555555556556656656666566556655566556655555555555555555568befffffffffffffffffffffffffffffffffffffffffff;
10'd406:mariog=956'hfffffffffffffffffffffffedba98888888888765555555555566666666555555555555555544544444444444434333333333333333333459bdfffff745555555555555555555555655665666566666665666566665565556555555555555555569dfffffffffffffffffffffffffffffffffffffffffff;
10'd407:mariog=956'hffffffffffffffffffffec9988887777777777776544455555555666666665555555555555555445444444444443333344333333333334458bcfffffa45555555555555555555555555665665566566656665566656665556555555555555555668bfffffffffffffffffffffffffffffffffffffffffff;
10'd408:mariog=956'hffffffffffffffffffeb988878777777777666666554444455555555666556555555455555445444444444444434333343333333333333447acfffffd44555555555555555555555556555655665566566665666566655565556555555555555567adffffffffffffffffffffffffffffffffffffffffff;
10'd409:mariog=956'hffffffffffffffffea88888877777777776666666555544444555555556555555555545555554454444444444443333353333333333333446abffffff645555555555555555555555655555566556666666566655666566655555565555555555559bffffffffffffffffffffffffffffffffffffffffff;
10'd410:mariog=956'hfffffffffffffffb98888887777777667666666655555444444445555555555555555544555555444444444444443334433333333333343459befffff955555555555555555555555555655665566556655666556666666556555555555555556667aefffffffffffffffffffffffffffffffffffffffff;
10'd411:mariog=956'hfffffffffffffda888888778777777766666666555555544444444455555555555555555455544444444444444434333433333333333334458adfffffc555555555555555555555555555556556656665566666666666555555555565566566666779cfffffffffffffffffffffffffffffffffffffffff;
10'd412:mariog=956'hffffffffffffc98888888777777777766666666655555544444444445555555555555555544554444444444444443434433333333333333457acffffff745555555555555555555655555665566556555666566666655556666666555555555667778beffffffffffffffffffffffffffffffffffffffff;
10'd413:mariog=956'hfffffffffffb888888888777777777766666666665555554444444444455555555555555554454444444444444444333443333333333333446abffffffa45555555555555555555555555555665565566666666655566666666555555555555555667adffffffffffffffffffffffffffffffffffffffff;
10'd414:mariog=956'hffffffffffb8888888877777777777777666666666555555544444444444445555555555555444444444444444444334433433333333333445abefffffc555555555555555555555555565566556556666666655566666666655655555555555555569bffffffffffffffffffffffffffffffffffffffff;
10'd415:mariog=956'hfffffffffa888888887777777777777777666666655555555544444444444454555555555555444544444444444444344433333333333334458beffffff7455555555555555565555555556556655666666656666666666655555555555555455455558dfffffffffffffffffffffffffffffffffffffff;
10'd416:mariog=956'hffffffffb8888888777777777777777666666666655555555544444444444344445555555444544444444444444443444333333333333334447bdffffffa4555555555555555555555555655665666666656666666666666655555555555545444445558fffffffffffffffffffffffffffffffffffffff;
10'd417:mariog=956'hfffffffc888888888777777777777777666666666555555554544444444444334544455545554445444444444444343444333333333333334469cffffffc4555555555555555555555555556656666665666666666665665555555554554444444454445affffffffffffffffffffffffffffffffffffff;
10'd418:mariog=956'hffffffd8888888878777777777777777776666666665555555444444444444443344444455445544444444444443433433343333333333334446afffffff65555555555555555555555555665666665566666666666566555555554554444444444343455bfffffffffffffffffffffffffffffffffffff;
10'd419:mariog=956'hffffff988888877777777877777777777777766666555555555444444444444443334444445544444444444444444434333333333333333344457cffffff855555555555555555555555565566666666666666666565555555554444444444333334334447dffffffffffffffffffffffffffffffffffff;
10'd420:mariog=956'hfffffb8888887777777877777777777777777776665555555554444444444444444334444444544444444444444344444434333333333334545569efffffa555555555555555555555565566666566666666666565555555544444444333323323323333359efffffffffffffffffffffffffffffffffff;
10'd421:mariog=956'hffffe98888777777777777788788878777777666666555555554444444444444444433444444444444444444444433444344443333333454444558bfffffc555555555555555555655555666656666666666656655555554444333322233344445566778889acefffffffffffffffffffffffffffffffff;
10'd422:mariog=956'hffffb88887777777777778888888888877777777666555555554444444444444444443334444444444444444444444343333333334444444444458bdffffe65555555555555555655655666656666666666555555555544443222233444455556666777788888899bdfffffffffffffffffffffffffffff;
10'd423:mariog=956'hfffe988777777777777788888888888888777777666665555554444444444444444444433344444444444444444444555444444444444443443448bcffffe65556555555555556556556665666666666666655555554443212334554455555566666677777777777879adffffffffffffffffffffffffff;
10'd424:mariog=956'hfffb877777777777777788888889988888887777666665555554444444444444444444443333444444444444444444454444444434334333333359bbfffff85555555555555555565665666666666666556555544433222345555555555566666666666777667777777778befffffffffffffffffffffff;
10'd425:mariog=956'hfff977777777777777778888899998988888777766665555555444444444444444444444433333344444444444444444444444343333333333346abbfffff7555555555555555565665666666666666555555444322234555555555555566666666666666666677777777778bffffffffffffffffffffff;
10'd426:mariog=956'hffd877777777777777778788899999889888787667665555555444444444444444444444444332333443343444443434544443333333333333347bacfffff755555555555555665655666666666665555555443223455555555555555666666666666666676776666776777779dffffffffffffffffffff;
10'd427:mariog=956'hffb77777777777777777878889999989988888777665555555554444444444444444444444433332333333333333334344333333333333333346abadffffd6555565555555555565666666666665555555443224555555555555556666666666666666777677776666777667777aeffffffffffffffffff;
10'd428:mariog=956'hff97777777777777777777889899999998888777766655555555444444444444444444444444333322233333333333334333333333233333345abbbeffffa555556555555555556766666666665555554432245555555555555556666666666666666676667666776666666777779dfffffffffffffffff;
10'd429:mariog=956'hfd87777777777777777788788888998988887777766655555554444444444444444444444444434443222233333333333333222222233333556abacfffff75555566556565665676666666565555555432245555555555555555556666666666666666666666677666666666776777cffffffffffffffff;
10'd430:mariog=956'hfc777777766666777777788888899988888887777666555555544444444444444444444444444444444322223222222322222222323334455558bbfffffd555555665656565566666666655555555433245555555555555555566666666666666666666667777777666666666676777afffffffffffffff;
10'd431:mariog=956'hfa777777666666666677778888888888888777777666555555544444444444444444444444444444444433222222233323233333333444444557acfffffb5555556655555566666666655555555443245555555555555555566666666666666666777777777777777676666666766677affffffffffffff;
10'd432:mariog=956'hf9777666666666667667778778888888878777776666555555544444444444444444444444444444444444432222223323333333333333444457abfffff8555566555665566666656655555545432245555555555555665566666666666666677777777777777777777766666666666779effffffffffff;
10'd433:mariog=956'hf87766666666666666667777888888888877777666655555555444444444444444444444444444444444444443322222233333333333334444569befffb65555556665556666666665555554542235555555555555555566666666666777777777777777777777777777766666666666779efffffffffff;
10'd434:mariog=956'he86666666666666666666777787788888877777666555555554444444444444443444444444444444444444444433333333333333333334444569bdfff756666656555666666656555555544322455555555555555566666666666777777777777777777777777777776766666666666677afffffffffff;
10'd435:mariog=956'hd76666666666666666666777777777777777776666555555555444444444443444444444444444444444444444434433333333333333344444559bcffc5566656655565666665555555544431355555555555555555566666666677777777777777777777777777777677666666666666677affffffffff;
10'd436:mariog=956'hd76666666666666666666666777777777777766666655555555444444444444444444444444344443344434443443444333333333333334444459bcffa55666655566666656565555554432135555555555556555666666666667777777777777777777777777777777666666666666666678bfffffffff;
10'd437:mariog=956'hc76666666666666666666666677777776766666665555555554444444444444444434443434444444444444444443344433333333333333444469bcff9566666656666665555555555443114555555555555555556666666667777777777777777777777777777777776666666666666666678cffffffff;
10'd438:mariog=956'hc7666666666666666666666666676666666666665655555555444444444444444434344343444434434444443444333333333333333333344446abcff96666565566666555555554543312455555555555555566666666666677777777777777777777777777777777666666666666666666679dfffffff;
10'd439:mariog=956'hc7666666666566665666666666666666666656655555555554444444444444444434334344433434333433333343333333333333333333344447abcffb6666666666555555555444432135555555555555556666666666677777777777777777777777777777777776666666666666666666668aeffffff;
10'd440:mariog=956'hd7666666666555555555556666666666666665565555555555444444444444444434344434334443333333333333333333333333333333344458badffd76666666555555555544433113555555555555555666666666666777777777777777777777777777777777766666666666666666666679cffffff;
10'd441:mariog=956'hd7666655655555555555555666666566666555555555555444444444444444444443334433343433333333333333333333333333333333344459badfff86666576555555544444321145555555555555556666666666667777777788888788777777777777777777777666666666666666666667aefffff;
10'd442:mariog=956'he766655555555555555555555566556655555555555555544444444444444444343334333334333433333333333333333333333333333344445abaefffb65555665555544444321024555555565655665556666666676777777788888888788777777777777777777676666666666666666666668cfffff;
10'd443:mariog=956'hf866555555555555555555555555565555555555555544444444444444444444333333333333333333333333333333333333333333333344447bbbfffff95555664545444443211355555555555566565566666666777777778878888888888787777777777777777666666666666666666666667adffff;
10'd444:mariog=956'hf965555555555555555555555555555555555555554444455444444444444443433333333333333333333333333333333333333333333334458bacffffff75554554444433311145555565555666566666666666666777777788888888888888777777777777777766666666666666666656666679bffff;
10'd445:mariog=956'hfa6555555555555555555555555555555555555554444444444444444444444444333333333333333333333333333333333333333333334446abbdffffffd6544554434321112455555555555555566566666666667777778888888888888888777777777777776766666666666666666665666668befff;
10'd446:mariog=956'hfc6555555555555555555555555555555555555555444444544444444444444433333333333333333333333333333333333333333333334458bbbeffffffd7555355332222235555555555565565665666666666677777888888888888888888777777777777766666666666666666666665555667acfff;
10'd447:mariog=956'hfd755555555555555555555555555555555555554444444444444444444444433333333333333333333333333333333333333333333334447abacfffffffc75544443333334555555665665566666556666666666777788898889999999888887777777776666666666666666666666665555566669bfff;
10'd448:mariog=956'hff85555555544445555555555555555555555554444444444444444444444333333333333333333333333333333333333333333333333446abbbefffffffc76544444444455566655666666666665566666666667777888989889999999898887777777766666666666666666666666555555556668adff;
10'd449:mariog=956'hffb5555555444444444445455555555555555554444444444444444444443333333333333333333333333333333333333333333333334469bbadffffffffc76655444455666666566666566556666665666666667777788889989899998888877777676776666666666666666666665555555555667acff;
10'd450:mariog=956'hfff755555444444444444444445455544445544444444444444444444433433333333333333333333333333333333333333333333345567ababfffffffffd766665556665666666666666666666566666666666677788888888998989988887777777776666666666666666665666555555555555679bef;
10'd451:mariog=956'hfffb65554444444444444444444444444444444444444444444444433333333333333333333333333333333333333333333333344555568abbffffffffffd766665556555666666666666666666555566666666667788888888899888888787777776666666666666666666655565555555555555669bdf;
10'd452:mariog=956'hffff85554444444444444444444444444444444444444444444444333333333333333333333333333333333333333333333444555555678abcffffffffffe766665555555566666666666666666555556666666677778788889998888887777777766666666666666666666655555555555555555568bcf;
10'd453:mariog=956'hffffe7555444444444444444444444444444444444444444444333333333333333333333333333333333333333333444545544455666678abcfffffffffff966565555655666666666665566666565665666666766677888888888888877777766666666666666666665555555555555555555555568bcf;
10'd454:mariog=956'hfffffd655444444444444444444444434444444444343343333333333333333333333333333333333333333344455444445555566666778abcfffffffffffa66655555556666666666665566666556565666666677677888888888888877777776666666666666666665555555555555555555555557abf;
10'd455:mariog=956'hffffffd7554444444443344444433344433433333333333333333333333333333333333333333333333334544444445555566666666668abacfffffffffffc66655555555556666666666666666566565566666667777777778887777777776666666666666666665565555555555555555555555557abe;
10'd456:mariog=956'hfffffffe8654444444433333343333333333333333333333333333333333333333333333333333333445554455555566666666666678abbbacfffffffffffe76655555556556666666666665555666655556666666767777777777777777777666666666666666655555555555555555555555555557abe;
10'd457:mariog=956'hffffffffa7655444433333333333333333333333333333333333333333333333333333333333434455555455556666666666666789abbbbabfffffffffffff96655555555555666666666656556565555556666666667677777777777766776666666666666655555555555555555555555555555557abe;
10'd458:mariog=956'hffffffffb976565443333333333333333333333333333333333333333333333333333333333345555555455666666666666789abbbbbaabdffffffffffffffc6655555555556666666666655556655555555556666666777777667777666666666666666555555555555555555555555555444455557abd;
10'd459:mariog=956'hfffffffebaa98655554433333333333333333333333333333333333333333333333333334455545567754456666667789abbbbbbaaabdefffffffffffffffff7665555555555666666666655555555555555555566666666666666776666666666655555555555555555555555555555444444455557bbd;
10'd460:mariog=956'hfffffffebaaaa99765555443333333333333333333333333333333333333333333333444555555668bba9766789aaabbbbbaaabbcdfffffffffffffffffffffa655555555555666666555555555555555555555656666666666666666666666666555555555555555555555555555544444444445557bbd;
10'd461:mariog=956'hfffffffebaaaaaaaa987654444333333333333333333322222333333333333333344545555566668bbbabbabbbbbbaaaaabcdefffffffffffffffffffffffffe765555555556666665555555555555555555555555666666666666666666656666655555555555555555555555555444444444445558bbe;
10'd462:mariog=956'hffffffffbabbbbaaaaaaa9987655443333333322222222232332333333333444445455556666679bbbadffdbaabbbcdeffffffffffffffffffffffffffffffffc65555555565666665555555555555555555555555566566656666666666655555555555555555555555555555544444444444445568bbe;
10'd463:mariog=956'hffffffffebabbbbbbaaaaaaaa9998776554444433333333333333333444444455555566666667abbbbdffffffefffffffffffffffffffffffffffffffffffffff95555555565666666655555555555555555555555555655666655655555555555555555555555555555555555544444444444445569bbe;
10'd464:mariog=956'hffffffffffbaabbbbbbbbbaaaaaaaa9999877665544444444444445455555555566666666668bbbabeffffffffffffffffffffffffffffffffffffffffffffffff8555555555666666655555555555555555555555555555565555555555555555555555555555555555555445444444444444445569bbf;
10'd465:mariog=956'hffffffffffebaaaaabbbbbbbbbaaaaaaaa9999998887665555555555556666666666666679bbbbabffffffffffffffffffffffffffffffffffffffffffffffffffe86555555566666655555555555555555555555555555555655555555555555555555555555555555544444444444444444444556abbf;
10'd466:mariog=956'hffffffffffffcbaaaaaabbbbbbbbaaaaaaaaa99999999988876666666666666666666679abbbabdffffffffffffffffffffffffffffffffffffffffffffffffffff97655555566666655555555555555555555555555555555555555555555555555555555555554544444444444444444444444557abcf;
10'd467:mariog=956'hffffffffffffffdbaaaa9aaabbbbaaaaaaaaaaa999999999998887766666666666679abbbbaacffffffffffffffffffffffffffffffffffffffffffffffffffffffb7666555566666655555555555555555555555555555555555555555555555555555555554445444444444444444444444444558bacf;
10'd468:mariog=956'hfffffffffffffffffdbbaaaa99aaaaaaaaaaaaaaa9999999998888887766667789bbbbbaabdffffffffffffffffffffffffffffffffffffffffffffffffffffffffba866666566666655555555555555555555555555555555555555555555555555555554444444444444444444444444444444569badf;
10'd469:mariog=956'hffffffffffffffffffffdcbbaaaaa999999999999999999988888877777889abbbbbaabceffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbaa9755666666665555555555555555555555555555555555555555555555555555555444444444444444444444444444444556abbef;
10'd470:mariog=956'hfffffffffffffffffffffffedcbaaabbbaaaa9999988888888888999aabbbbbbaaabdefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdaaaa86556666666555555555555555555555555555555555555555554444445555444444444444444444444444444444444557abbff;
10'd471:mariog=956'hffffffffffffffffffffffffffffedccbbbaaabbbbbbbbbbbbbbbbbbbaaaabbcdeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcaaaa9766677666555555555555555555555555555555555555555555555444444444444444444444444444443343344444559bacff;
10'd472:mariog=956'hfffffffffffffffffffffffffffffffffffeddcccbbbbbbbbbbbbbbbccddeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcaaaaa8666676655555555555555555555555555555455545554555555444444444444444444444444444433333334444556abadff;
10'd473:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc9aaaa976657665555555555555555554444444555555555444444444444444444444444444444443443333333344444558bbbfff;
10'd474:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdaaaaaa864486655555555555545454444455555555555444444444444444444444444444444433333333333334444456abacfff;
10'd475:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffebaa9aa84478655555544554544444444445445555554444444444444444444444444444443333333333333333444458bbbdfff;
10'd476:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecaaaa646976555555444444444444444444444544444444444444444444444444443333333333333333333444457abacffff;
10'd477:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbaaaba8765554444444444444444444444444444444444444444444444443333333333333333333333344446abbbeffff;
10'd478:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbaaa876554444444444444444444444444444444444444444444333333333333333333333333333444458bbacfffff;
10'd479:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecaa8665544444444444444444444444444444444444434433333333333333333333333333333344458bbabffffff;
10'd480:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbaa86655444444444444444444444444444444443333333333333333333333333333333333444458bbbbeffffff;
10'd481:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeaa9866554444444444433333444444434333333333333333333333333333333333333333344468bbbadfffffff;
10'd482:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcaaa976654444444443333333333333333333333333333333333333333333333333333444457abbbadffffffff;
10'd483:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffbaaa9976554443333333333333333333333333333333333333333333333333333334444567abbabdfffffffff;
10'd484:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeaaaa998755544433333333333333333333333333333333333333333333333333444556667ababeffffffffff;
10'd485:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdaaaaa9997655544333333333333333333333333333333333333333333333344555555678abaefffffffffff;
10'd486:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdaaaaaa99987655544333333333333333333333333333333333333344445555555566778abaefffffffffff;
10'd487:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd9aaaaaa999987654444433333333333233333333333333344445555555555566667778abaefffffffffff;
10'd488:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdaaaaaaaaaa99998765544444444433333344444445455555554455555566666777779abaefffffffffff;
10'd489:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffea9aaaaaaaaaaa999988765544444544544445544455555555555666666667777778abbbffffffffffff;
10'd490:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb99aaaaaaaaaaaaa9999998776555555555555555556666666666666777777778abbacffffffffffff;
10'd491:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda99aaaaaaaaaaaaaaaa9999999988766666666666666666666667777777789bbbabfffffffffffff;
10'd492:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcba99aaaaaaaaaaaaaaaaaaaa999999988777666666667667777776778abbbbabffffffffffffff;
10'd493:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecaaa99aaaaaaaaaaaaaaaaaa99999999999888777677766666678aabbbaabdfffffffffffffff;
10'd494:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdbaaa99999aaaaaaaaaaaaaa99999999999999877667789abbbbbaaabdfffffffffffffffff;
10'd495:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbbaaaa99999999999999999999988888888899aabbbbbaaabcdffffffffffffffffffff;
10'd496:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedcbaabaaaa99998888888999999aaaabbbbbbbaaaabcdefffffffffffffffffffffff;
10'd497:mariog=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdccbbaabbbbbbbbbbbbbbbbbbaaaaaabbccdeffffffffffffffffffffffffffff;
10'd498:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeddcbbbbbbbbbbbbbbcccddeefffffffffffffffffffffffffffffffffff;
10'd499:mariog=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;


	endcase
	case((y_cnt-move_y))
 10'd0:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedcba9888778899abcdefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd1:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeca86554433333333333333444568acefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd2:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffca75443333333333333333333333333333467adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd3:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda7443333333332222222222222222223333333333347adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd4:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffea7544333333222222222222222222222222222223333333346aeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd5:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd8543333333222222222222222222222222222222222222333333347bffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd6:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc643333333222222222222222222222211212112122222222222233333338dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd7:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffc7443333322222222222222222222222212111111111112222222222223333346cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd8:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffd84333333222222222222222222222222221211111111111111122222222233333335bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd9:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffff944333322222222222222222222222222221111111111111111111122222222223333335afffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd10:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffc743333222222211111122222222222222222121111111111111111111111222222223333335bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd11:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffff9543332222100246777642001222222222121111111111111111111111111111222222223333336cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd12:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffe843333221126aefffffffffeb521122212221111111111111111111111111111111212222223333337dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd13:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffe7433322214aeffeddddddedefffe92112211121111111111111111111111111111111122222223333335affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd14:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffe643322213cffedeeffffffbeeddffff81112121111111111111111111111111111111111122222223333336dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd15:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffc63332212affedfffffffffb39fffddeffe30111111111111111111111111111111111111111122222223333348fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd16:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffc64332214efeeffffffffffd645effffdefff50111111111111111111111111111111111111111122222223333346dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd17:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffd54332218ffeffffffffffff75538fffffedeff60111111111111111111111111111111111111111112222222233334affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd18:mariob=956'hffffffffffffffffffffffffffffffffffffffffffd7433221afedffffffffffffb55445dffffffdeff501111111111111111111111111111111111111111112222222333437effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd19:mariob=956'hffffffffffffffffffffffffffffffffffffffffff84332219fee6bffffffffffd6554448fffffffdefe301111111111111111111111111111111111111111112222222333345cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd20:mariob=956'hfffffffffffffffffffffffffffffffffffffffff94332219fefc549fffffffff75544444bfffffffdffc111111111111111111111111111111111111111111111222222333344affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd21:mariob=956'hffffffffffffffffffffffffffffffffffffffffb4433217feff95549fffffffa555444444dfffffffeff70111111111111111111111111111111111111111111112222222333447effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd22:mariob=956'hfffffffffffffffffffffffffffffffffffffffd6433213feffd655548fffffd65554444437fffffffeffd11111111111111111111111110110111111111111111111222222333446efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd23:mariob=956'hfffffffffffffffffffffffffffffffffffffff7433222cfeffc5455547ffff855554444444afffffffeff601111111111111111101111111101111111111111111111122222333345cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd24:mariob=956'hffffffffffffffffffffffffffffffffffffffa4332217fefff954555557efb5554444444445dffffffeffb111111111111111111111011100101111111111111111111222222333344afffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd25:mariob=956'hfffffffffffffffffffffffffffffffffffffe5432222deffff7545555547e755544434444448fffffffffe3011111111111110111010110101011011111111111111111222222233344affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd26:mariob=956'hfffffffffffffffffffffffffffffffffffff84332218fffffc54445555555555544443444443bffffffeff701111111111111101000001000001010111111111111111111222222333448fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd27:mariob=956'hffffffffffffffffffffffffffffffffffffb5332212efffff954445555455554543c934444444cffffffefa011111111110101110100100000000011110111111111111111122222333448ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd28:mariob=956'hffffffffffffffffffffffffffffffffffff74332215fefffe644444545555545536fd434444446ffffffffb1011110101010111000100000000000000100111111111111111222222333448fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd29:mariob=956'hfffffffffffffffffffffffffffffffffffb4432211afffffc54443345545554443cff8344444437fffffefd10111110101010001010000001000000100110111111111111111122222333447ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd30:mariob=956'hfffffffffffffffffffffffffffffffffff74322213efffffb54443964545554436fffd344444444dffffeed201000110101011000010100000000000000101101111111111111122222333447fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd31:mariob=956'hffffffffffffffffffffffffffffffffffc44322216ffffff954443cf644555443bffff5344444445dfffeed2000101000000001000010000000000000000001111111111111111112222333448ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd32:mariob=956'hffffffffffffffffffffffffffffffffff743322209ffffff744434dff63455435fffffc3444444437fffffd30100000000000000000000000000000000001000101111111111111122222233447fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd33:mariob=956'hfffffffffffffffffffffffffffffffffc54322211bfffffd644434dfff534543affffff7344444444affffd200000000000000000000000000000000000000001001111111111111122222333448ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd34:mariob=956'hfffffffffffffffffffffffffffffffff943322211cfffffb544434efffe53444effffffc3344434444cfffc1000000000000000000000000000000000000000001010111111111111112222333449fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd35:mariob=956'hffffffffffffffffffffffffffffffffe643222212efffff8444435efffff6338ffffffff63344444445dfeb10000000000000000000000000000000000000000010010111111111111122222333459ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd36:mariob=956'hffffffffffffffffffffffffffffffffb543222113efffff7444435fffffff53dffffffffd33434444438fe900000000000000000000000000000000000000000000011111111111111111222233445bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd37:mariob=956'hffffffffffffffffffffffffffffffff8433222113eefffc5544436fffffffeaffffffffff7334443433bfe7000000000000000000000000000000000000000000000010111111111111112222233446cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd38:mariob=956'hfffffffffffffffffffffffffffffffe6433221112effffc5444437fffffffffffffffffffe43443432afed40000000000000000000000000000000000000000000000010011111111111111222233446cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd39:mariob=956'hfffffffffffffffffffffffffffffffc5432221112dffffb5444428ffffffffffffffffffff92333427efeb200000000000000000000000000000000000000000000000100111111111111111222233447effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd40:mariob=956'hfffffffffffffffffffffffffffffffa4332221111cffff84444428ffffffffffffffffffffe533424defe80000000000000000000000000000000000000000000000000000111111111111111222233458ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd41:mariob=956'hfffffffffffffffffffffffffffffff743322211109efff84444429fffffffffffffffffffefb2324cdfec400000000000000000000000000000000000000000000000000000110111111111111222233459fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd42:mariob=956'hffffffffffffffffffffffffffffffd643322111107fffe6444442affffffffffffffeeeeeeee622addfda100000000000000000000000000000000000000000000000000000011111111111111122233345affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd43:mariob=956'hffffffffffffffffffffffffffffffc543222111103effd5444442afffffffffffefeffeeeeeeb27ddfec60000000000000000000000000000000000000000000000000000000001111111111111222233446cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd44:mariob=956'hffffffffffffffffffffffffffffffa543222111111affc5444442bffffffeeeeeeeeeeeeedded9ccefc9100000000000000000000000000000000000000000000000000000000101111111111111122233447dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd45:mariob=956'hffffffffffffffffffffffffffffff84432221111105ffb4444443bffffeefeeeeeeeeeeddddeeddeedb50000000000000000000000000000000000000000000000000000000000011111111111111222233448efffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd46:mariob=956'hffffffffffffffffffffffffffffff74332221111101cfc4344433bfeeeeeeeeeededdddddeeeeeeedb7000000000000000000000000000000000000000000000000000000000000101111111111111222233459fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd47:mariob=956'hfffffffffffffffffffffffffffffe643322211111105ffe843432bfeeeeeeddddddeefeeeedddddcb81000000000000000000000000000000000000000000000000000000000000000011111111111122223345cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd48:mariob=956'hfffffffffffffffffffffffffffffd643322111111100affec6333beeeeddddddeeeedddccba975543221110000000000000000000000000000000000000000000000000000000000001011111111111222223347dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd49:mariob=956'hfffffffffffffffffffffffffffffc5433221111111001cffeea419eedddcdffedddcb9754333334333322111111111110000000000000000000000000000000000000000000000000010111111111111222223359effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd50:mariob=956'hfffffffffffffffffffffffffffffb54332211111111102dffeee99ddddeeedcca75444444444443433332221111111111111100000000000000000000000000000000000000000000001101111111111122222345affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd51:mariob=956'hfffffffffffffffffffffffffffffa543222111111000003cefedddcdefedb8654445544444443333333322222111111111111111111000000000000000000000000000000000000000000111111111111122223347dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd52:mariob=956'hfffffffffffffffffffffffffffff95432221111111100002beffdcdfec86445544444444444433333333322222221121111111111111110000000000000000000000000000000000000000111111111111122223348dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd53:mariob=956'hfffffffffffffffffffffffffffff8443222111111100000007cdefe9644455555545444433333333333332222222222221111221111111111000000000000000000000000000000000000011111111111112222233569effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd54:mariob=956'hfffffffffffffffffffffffffffff844322211111110000000039b85445555444333332222222222222222222222222222222222221111111111000000000000000000000000000000000000111111111111122222345569effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd55:mariob=956'hfffffffffffffffffffffffffffff8443221111111000000000134444443333322222222111211111111111111112222222222222222211111111110000000000000000000000000000000000111111111111122222355555bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd56:mariob=956'hfffffffffffffffffffffffffffff744322211111100000013444433333222211111100010000000000000000000000011111222222222222222111110000000000000000000000000000000001111111111111222234545557dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd57:mariob=956'hfffffffffffffffffffffffffffff7443222111111100023444332221111100000000000000001001001000000000001000000111122222222222211111000000000000000000000000000000011111111111112222235444455cffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd58:mariob=956'hfffffffffffffffffffffffffffff74432221111100134433221111000000000000000100110011011010010010000000001000000001122222222222211100000000000000000000000000000111111111111112222344444445afffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd59:mariob=956'hffffffffffffffffffffffffffffe7443222111113443322110100000000000011111111111111111111111111111111000000000000000011222222222221100000000000000000000000000011111111111111122223433444459ffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd60:mariob=956'hffffffffffffffffffffffffffffe74432211134432111100000000001111111111111111111111111111111111111111111110100000000000012222222222110000000000000000000000000011111111111111122223333344459fffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd61:mariob=956'hfffffffffffffffffffffffffffff744322345421111100000000111111111111111111111111111111111111111011001111111111000000000000122222222211000000000000000000000000010111111111111122223333334459ffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd62:mariob=956'hfffffffffffffffffffffffffffff743345421000100000011111111111111111111111111111111111111111111110001000101111111111001010000122222222210000000000000000000000011111111111111112222223333445afffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd63:mariob=956'hfffffffffffffffffffffffffffff7555411000010001111111111111111111111111111111111111111111111100000000000001111101111100001100012222222111000000000000000000000011111111111111112222222333446cffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd64:mariob=956'hfffffffffffffffffffffffffffff84310100001111222111111111111111111111111111111111111111111000000000000000000000011111111100011001122222221000000000000000000000011111111111111122222222333448dfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd65:mariob=956'hfffffffffffffffffffffffffffd7211001100112222211111111111111111111111111111111111112222233333333321000000000000000000011110001000112222221100000000000000000000111111111111111111222222333459effffffffffffffffffffffffffffffffffffffffffffffffff;
10'd66:mariob=956'hffffffffffffffffffffffffff931011001112222221111111111111111111111111111111122333444444444444443310000000000000000011100111110010011122222100000000000000000000011111111111111111122222233447cffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd67:mariob=956'hffffffffffffffffffffffffc40000111122222222222111111111111111111111111123344444444444444444444420000000000000000000134433211111111111122222210000000000000000001011111111111111111122222233458efffffffffffffffffffffffffffffffffffffffffffffffff;
10'd68:mariob=956'hfffffffffffffffffffffff9110010112222222222111111111111111111111111223444444444444444555555444200000000000000000000023344443321111111111222211000000000000000001111111111111111111112222223346bfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd69:mariob=956'hfffffffffffffffffffffe71110011222222222222211111111100000111111133444444444444555555555555443000000000000000000000003344444443321111111122221100000000000000001011111111111111111111222223345adffffffffffffffffffffffffffffffffffffffffffffffff;
10'd70:mariob=956'hffffffffffffffffffffe3110011223322222222221111111000000000011244444444444555555555555555554300000000000000000000000013444444444433111111122222000000000000000001111111111111111111111222223348befffffffffffffffffffffffffffffffffffffffffffffff;
10'd71:mariob=956'hfffffffffffffffffffd41101122222222222222111111110000000001234444444445555555555555555555554100000000000001111100000002444444444444331111111222110000000000000000011111111111111111111122223346adfffffffffffffffffffffffffffffffffffffffffffffff;
10'd72:mariob=956'hffffffffffffffffffd4001012223222222222221111111111000000234444444455555555555555555555555520000001111111111110000000014445544444444432111111122110000000000000001011111111111111111111222233359bfffffffffffffffffffffffffffffffffffffffffffffff;
10'd73:mariob=956'hfffffffffffffffffe31111222322222222222211111110000000023444444455555555555555555555555555410011111111111111111111100003555555554444444421111111111000000000000011111111111111111111111122223358beffffffffffffffffffffffffffffffffffffffffffffff;
10'd74:mariob=956'hfffffffffffffffff610112222222222222222121111110000001334444555555555555555555555555666555200111111111110101000111111002555555555555444443211111111000000000000011111111111111111111111112223347adffffffffffffffffffffffffffffffffffffffffffffff;
10'd75:mariob=956'hffffffffffffffff9111122222222222222222211111000000122234444555555555555555555556566666554101111111110011223332110011101455555555555555544432100001000000000000001111111111111111111111112223346acffffffffffffffffffffffffffffffffffffffffffffff;
10'd76:mariob=956'hfffffffffffffffc2111222222323222222222211111100001000001344555555555555556666666666666653011111110012445555555554310110355565555555555555554420000000000100000011111111111111111111111111222346abffffffffffffffffffffffffffffffffffffffffffffff;
10'd77:mariob=956'hfffffffffffffff611122222222222222222221111110000000000000245555555556565666666666666666520111111123455566666666666531002566666666566556656555420000000000101000111011111111111111111111112223459befffffffffffffffffffffffffffffffffffffffffffff;
10'd78:mariob=956'hffffffffffffffd211122222222222222222221111000000000000000024555555566566666666666666666511111101355666666666666666666302566666666666666666666530000000000011011110111111111111111111111112223359bdfffffffffffffffffffffffffffffffffffffffffffff;
10'd79:mariob=956'hffffffffffffff7111222222222222222222221111000010000011000002455566666666666666666666666411111025666666666666666666666641566666666666666666666651000000000011111101111111111111111111111112223359bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd80:mariob=956'hfffffffffffffe4111222222222222222222211111000100000111100000355566666666666666666666666301111356666666666666666666666665666666666666666777777662000000000000011111111111111111111111111112223359bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd81:mariob=956'hfffffffffffffd4212222222222222222222221110001100011111110000145666666666666666666666666301103666666766777677777666666667766666666677777777777774000000000100001111111111111111111111111112223359bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd82:mariob=956'hfffffffffffffb3112222222222222222222211110002001111111110010025666666666666666666666666211136767777777777777777777777777777777777777777777777775000000000111000011111111110111111111111112223359bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd83:mariob=956'hfffffffffffffb2122222222222222222222211100012011111111111101004666666666666666666666666211367777777777777777777777777777777777777777777777777776000000000111110011111111111101110111111112223359bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd84:mariob=956'hfffffffffffffc312222222222222222222211111002201111111111111110356666666666666666666666620257777777777777777777777777777777777777777777777777777610000000001112100111111000000000001111111122335abcfffffffffffffffffffffffffffffffffffffffffffff;
10'd85:mariob=956'hfffffffffffffc322222222222222222222111110003101111222222221110156666666666666666666667621567777776666666667777777777777777777777777777777777777720000000001122220011000000000000000011111222335abcfffffffffffffffffffffffffffffffffffffffffffff;
10'd86:mariob=956'hfffffffffffffd422222222222222222222111000014111122222222222111046666666666666666667677623677777666666777666677777777777777777777777777777777777720000000001122222000000000000000100000111222346abcfffffffffffffffffffffffffffffffffffffffffffff;
10'd87:mariob=956'hffffffffffffff7112222222222222222221111000240112223444443322210266666666666666666777777467777776679bbcccca8666777777777777777777777777777777777720000000001122222200000000035678888764101222347aacfffffffffffffffffffffffffffffffffffffffffffff;
10'd88:mariob=956'hffffffffffffffb212222221222222222221110000341112345555555554320156666666666667777777777777777667accccccccccc96677888888888888888888788878888877720000000001122222210000015788888888899973122348badfffffffffffffffffffffffffffffffffffffffffffff;
10'd89:mariob=956'hfffffffffffffff51222222222222222222111000044111455666666666543104666666667777777888888888777769bcccccdcdccccca778888999998888888888888888888877730000000000122222220000278888888888888899612348bbdfffffffffffffffffffffffffffffffffffffffffffff;
10'd90:mariob=956'hfffffffffffffffb212221221222112221111100004411356666666666666531376666777777888888888888887769ccddddddddddddddb77889999999999998899888888888887730000000000122222210004788888888888888888a72359bbefffffffffffffffffffffffffffffffffffffffffffff;
10'd91:mariob=956'hffffffffffffffff92222221111212112111100000441256666666777777665326777777788888888888888888768cdddddddddddddddddc778999999999999999899998888888873000000000012222221004789999999888888888889836abbffffffffffffffffffffffffffffffffffffffffffffff;
10'd92:mariob=956'hfffffffffffffffff622221121112211111111000055146666667777777777664677778888888888888888888777bddddeedeeeeeeddddddb78899999999999999998988888888873000000000112222321027899999988888888888888987aacffffffffffffffffffffffffffffffffffffffffffffff;
10'd93:mariob=956'hffffffffffffffffff6221211211111111111110005526666667777777777777667788888888888888888888877acddddeeeeeedccbccccdd9789999999999999999989898888887300000000011222232016899999988888888888888889abadffffffffffffffffffffffffffffffffffffffffffffff;
10'd94:mariob=956'hfffffffffffffffffff832222111111111111110015666667777777766677777778888888888888888888888878bdddeeeeeedbbcccdddcbcc878999999999999999999999888887200000000011222332048999999888888888888888888abaeffffffffffffffffffffffffffffffffffffffffffffff;
10'd95:mariob=956'hffffffffffffffffffffb5212221111111111111105777777777766669aba977788888888888888888888888779cddeeeeeecbccdddddddcbca789999999999999999999998888861001000001122222321689999888887777777788888889abfffffffffffffffffffffffffffffffffffffffffffffff;
10'd96:mariob=956'hfffffffffffffffffffffd9522222222211111111057777777777655bddcddc978888888888888888888888877bddeeeeeecacdddddddddddbc789999999999999999999999888850010000111122223323799998888776666666677888888abeffffffffffffffffffffffffffffffffffffffffffffff;
10'd97:mariob=956'hffffffffffffffffffffffeca753322222222222216877777777655bdccddddda7888888888888888889988878bdeeeeeedacdddddddddccddc9789999999999999999999998887401111111111222223258999888877666666666677888889acffffffffffffffffffffffffffffffffffffffffffffff;
10'd98:mariob=956'hffffffffffffffffffffffffdbba977656677886317977777777649dddddddddea888888888888888899988879cddeeeeebbdddddddddcccddda789999999999999999999998886201111111112222233268988888776666666766667788888abefffffffffffffffffffffffffffffffffffffffffffff;
10'd99:mariob=956'hffffffffffffffffffffffffffecbbbbbbbbbbbb93798777777656cddddeeeedcb888888888888899999988879cddeeeedadddddeda9acddccdb7899999999999999999999888840110111111122223333788888877666777777777667888889bcfffffffffffffffffffffffffffffffffffffffffffff;
10'd100:mariob=956'hfffffffffffffffffffffffffffffeccbbbbbbbbc87a8777777649ddddddddbbbba8888888888888999999887adddeeeebbddddea543349dccdd8799999999999999999999988821111111111222222333788888776777788887777777788889abeffffffffffffffffffffffffffffffffffffffffffff;
10'd101:mariob=956'hffffffffffffffffffffffffffffffffffffffffffba887777764cdddddddcccddca888888888889999999887addddeeeacdddeb44344338dcde9789999999999999999999888711111100011222222334788888777778888888877777788888abdffffffffffffffffffffffffffffffffffffffffffff;
10'd102:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffb888777755dddddedcddddccc888888888889999999887bdddddedaddcdc434aed533bddda689999999999999999999988611111111111222222334788887777888888888888777788888abcffffffffffffffffffffffffffffffffffffffffffff;
10'd103:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffb888777757eedeedcdddddccc988888888889999999887bddddddcacccd8238fffa337dcdc6899999999999999999998885111111100112232223357888777778888888888888777888889bbffffffffffffffffffffffffffffffffffffffffffff;
10'd104:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffc988777759eeeeeddeddddcccb88888888889999999887bddddddbaccdd533afffc334bddb6899999999999999999998885111111000122321123467888777788888888888888877888889bbefffffffffffffffffffffffffffffffffffffffffff;
10'd105:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffd98888875aeeeedcddddc6477998888888899999999887bddddddbadcdb3336fff83328ddc6889999999999999999999885111111100112201223467888777777788888888888877788889aaefffffffffffffffffffffffffffffffffffffffffff;
10'd106:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffd98888876bddeeddeddb43dfc378888888899999999887bddddddbaccdb33337b833326ddd6889999999999999999999886111111000123001223567887777777778888888888887788889aadfffffffffffffffffffffffffffffffffffffffffff;
10'd107:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffe98888877cdddeddedc436fff458888888899999999887addddddabccdb333333333334cdd7789999999999999999999987101110001122001123567887776655566788888888887788889aacfffffffffffffffffffffffffffffffffffffffffff;
10'd108:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffea9998877dddddcddd9234ffc348888888899999999887addddddaaccdb333344444333bdd8789999999999999999999988200000001120011223577777665555555678888888887788889aacfffffffffffffffffffffffffffffffffffffffffff;
10'd109:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffa9998878dddddcddd623258423788888889999aa998879ddddddaaccdc333456776433bee8789999999999999999999999600000001100001223577776666666655557888888887788889aacfffffffffffffffffffffffffffffffffffffffffff;
10'd110:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffb9998878dedddceed43566677689888888999aaa998878cdddddb9ccdc434468aa8543aee9799999999999999999999998830000010001011223577776666667776666788888897888889bbcfffffffffffffffffffffffffffffffffffffffffff;
10'd111:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffc9999878dddedcdb999999999988899998999aaa999878bdcdddc9cbcd63459bdca743aeea799999999999999999999999883000000000001123677766666777888766688888898888889abcfffffffffffffffffffffffffffffffffffffffffff;
10'd112:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffca999888dedca988899888888888888889999aaa999887bdcdddc8bcce9246adeeb844beea899999999999999999999999888411000110011223677766667778888876678888998888889bacfffffffffffffffffffffffffffffffffffffffffff;
10'd113:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffda999887db989999999999999998888888899aaa998887adcccdd9cdcdb346adeec844dee9899999aaa999999999999999988873001110011223677766667788888877678888998888889bacfffffffffffffffffffffffffffffffffffffffffff;
10'd114:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffda999889989999999999999999999999888888999988878cccccdaadcde5369cddb747efd899aaaaaaa999999999999999999885001100011223677766677888888887678888998888889badfffffffffffffffffffffffffffffffffffffffffff;
10'd115:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffea9999a9999999999999999999999999998888899988887bccccdc9cddeb358abb963affb89aa99996389888889999999999988710111000122467776677888888888777888899898888abadfffffffffffffffffffffffffffffffffffffffffff;
10'd116:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffb99aa999999999999999999999999999998888899988879cccccd9bedef736888746ffe8899988972148888888999999999998830110000112477776678888888888777888899898888abaefffffffffffffffffffffffffffffffffffffffffff;
10'd117:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffcaaa99999999999999aa999999999999999998888998888bccccdb9eeeef8355535fff97888888712225988888989999999999961011000112477776678888888888777888999998889bbbefffffffffffffffffffffffffffffffffffffffffff;
10'd118:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffcbaa99999999999aaaaaaaaa9a9999999999999889998879cccccc9bfeeffc866afffc78888886222222788888889999999999983000000112577776778888888998777989999988889bbbffffffffffffffffffffffffffffffffffffffffffff;
10'd119:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffdaa9999999999aaaaaaaaaaaaaa999999999999988899887acccccc9dfffffffffffb7888889622222224888888899999999999970000001226777767888888899988789999aa98888abbcffffffffffffffffffffffffffffffffffffffffffff;
10'd120:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffba999999999aaaaaaaaaaaaaaaaaa99999999999988999888bcccccb9cffffffffe97888888512222222278888888899999999999500001123777776788888899999778999aa988888bbbdffffffffffffffffffffffffffffffffffffffffffff;
10'd121:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffcaa999999999aaaaaaaaaaaaaaaaaaa99999999999888999888bcccccb9ceffffea878888874122222222248888888889999999999820001125777777788888899998789999aa988889bbbeffffffffffffffffffffffffffffffffffffffffffff;
10'd122:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffeaaaa9999999aaaaaaaaaaaaaaaaaaaa999999999999888998888abccccc9accb9778888886212222222222378888888889999999999710111487777877888889999977999aaa998888ababfffffffffffffffffffffffffffffffffffffffffffff;
10'd123:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffbaa999999999aaaaaaaaaabbbbbaaaaaa999999999999888998888899aa99877778888886312222333222222688888888888999999999711258877778778888889997799aaaa9988889bbadfffffffffffffffffffffffffffffffffffffffffffff;
10'd124:mariob=956'hffffffffffffffffffffffffffffffffffffffffffdaaa9999999999aaaaaaaaaabbabaaaaaa9999999999998888987888888877888888888631222223333322222588888888888999999999974688877788888888889988899aaaa998888abbbefffffffffffffffffffffffffffffffffffffffffffff;
10'd125:mariob=956'hffffffffffffffffffffffffffffffffffffffffffcaa9999999999aaaaaaaaaaabbbaaaaaaaa99999999999888889888888888888888885212222222333332222247888888888888999999999888888778889888888888899999a9988888bbacffffffffffffffffffffffffffffffffffffffffffffff;
10'd126:mariob=956'hfffffffffffffffffffffffffffffffffffffffffebaa99999999999aaaaaaaaaaabaaaaaaaaa9999999999988888888888888888888632122222223333333222223788888888888899999999998888887888888888888888999999888889bbaeffffffffffffffffffffffffffffffffffffffffffffff;
10'd127:mariob=956'hfffffffffffffffffffffffffffffffffffffffffdaaa999999999999aaaaaaaaaaaaaaaaaaa9999999999998888888788888888874211222222223333333222222368888888888888999999999988888788888888888888889999888888ababfffffffffffffffffffffffffffffffffffffffffffffff;
10'd128:mariob=956'hfffffffffffffffffffffffffffffffffffffffffcaa9999999999999aaaaaaaaaaaaaaaaaaa999999999998888888878889876421122222222233333333322222236788888888888889999999999988878888888888888889999988888abbadfffffffffffffffffffffffffffffffffffffffffffffff;
10'd129:mariob=956'hfffffffffffffffffffffffffffffffffffffffffbaa99999999999999aaaaaaaaaaaaaaaaaa999999999998888888777764321222222222223333333333222222246788888888888889899999999988888888888888888889998888889bbacffffffffffffffffffffffffffffffffffffffffffffffff;
10'd130:mariob=956'hffffffffffffffffffffffffffffffffffffffffebaa99999999999999aaaaaaaaaaaaaaaaa999999999998888888874221122222222222223333333333322222124678888888888888889999999999888888888888888888998888888abbbeffffffffffffffffffffffffffffffffffffffffffffffff;
10'd131:mariob=956'hffffffffffffffffffffffffffffffffffffffffeaa9999999999999999aaaaaaaaaaaaaaa9999999999999888888773122222222222222333333333332222222236678888888888888889899999999888888888888888888888888889bbacfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd132:mariob=956'hffffffffffffffffffffffffffffffffffffffffeaa999999999999999999aaaaaaaaaaa99999999999999888888877312222222222222333333333332222222114667888888888888889899999999998888888888888888888888889bbbbefffffffffffffffffffffffffffffffffffffffffffffffff;
10'd133:mariob=956'hffffffffffffffffffffffffffffffffffffffffeaa99999999999999999999a9aaa99999999999999998888888887731222222222222333333333322222222122666788888888888888989999999999888888888888888888888878abbadffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd134:mariob=956'hffffffffffffffffffffffffffffffffffffffffeaa99999999999999999999999999999999999999999888888887762222222222222333333333222222222112466678888888888888888999999999988888888888888888888878abbacfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd135:mariob=956'hffffffffffffffffffffffffffffffffffffffffeaa9999999999999999999999999999999999999998888888888776222222222222333333332222222222111466667888888888888888889999999998878888888888888888878abbabefffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd136:mariob=956'hffffffffffffffffffffffffffffffffffffffffeba999999999999999999999999999999999999999888888888877512222222322333333332222222222111366667888888888888888888899999999877788888888888888878abbbaeffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd137:mariob=956'hfffffffffffffffffffffffffffffffffffffffffba99999999999999999999999999999999999998888888888877732223333333333333333222222211111366667788888888888888888889999999987677788888888877778abbbadfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd138:mariob=956'hfffffffffffffffffffffffffffffffffffffffffca9999999999999999999999999999999999988888888888877762233333333333333333222222111112466667788888888888888888888899999998656677777777777779abbbbdffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd139:mariob=956'hffffffffffffffffffffffffffffffffffffffffc9a99999999999999999999999999999999988888888888887777413333333333333333332222111111356666777888888888888888888888999999996556667777777778abbbaaefffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd140:mariob=956'hffffffffffffffffffffffffffffffffffffffff67b9999999999999999999999999999999888888888888888777622333333333333333333222222123566666777888888888888888888888899999aa963556666666778abbbbabeffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd141:mariob=956'hfffffffffffffffffffffffffffffffffffffffc34ba99999999999999999999999999988888888888888888777741333333333333333222222222235556666777888888888888888888888889999aaa9612356677778abbbbaadffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd142:mariob=956'hfffffffffffffffffffffffffffffffffffffff9329a99999999999999999999999989888888888888888877777612333233333333322222222222245566667788888888888888888888888889999aaa96111122223248bbaacefffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd143:mariob=956'hfffffffffffffffffffffffffffffffffffffff7325b99999999999999998988888888888888888888888777777312222222222222222222222222245666677888888888888888888888888889999aaa941111111112349bdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd144:mariob=956'hffffffffffffffffffffffffffffffffffffffe53327a9999999888888888888888888888888888888888777775112222222222222222222222212256667788888888888888888888888888889999aaa821111111112236bfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd145:mariob=956'hffffffffffffffffffffffffffffffffffffffe43323ba99998988888888888888888888888888888887777776212222222222222222222222211235678888888888888888888888888888889999aaaa6111111111112259dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd146:mariob=956'hffffffffffffffffffffffffffffffffffffffd433214a99988888888888888888888888888888888777777772012222222222222222222221111246678888888888888888888888888888889999aaaa3111111001111238befffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd147:mariob=956'hffffffffffffffffffffffffffffffffffffffd4332216a9988888888888888888888888888888777777777730122221112222222222222211112266688888888888888888888888888888889999aaa81001100000111238adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd148:mariob=956'hffffffffffffffffffffffffffffffffffffffd43322227b988888888888888888888888888887777777777401122221112222222222222111111466788888888888888888888888888888889999aab50111011010111248bbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd149:mariob=956'hfffffffffffffffffffffffffffffffffffffff622222226a9888888888888888888888878777777777777301122222111112222222221111111366778888888888888888888888888888888999aab910000010000011248bbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd150:mariob=956'hfffffffffffffffffffffffffffffffffffffff9322222326a988888888888888888888877777777777773011222222211112221112111111112667778888888888888888888888888888888999aab600000000000111249bbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd151:mariob=956'hfffffffffffffffffffffffffffffffffffffffe62222233239a9888888888888888777777777777777620111222222221111111111111111126667778888888888888888888888888888889999aba20010111110011226abbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd152:mariob=956'hffffffffffffffffffffffffffffffffffffffffe522223332159a8888888888777777777777777777400111221122221111111111111111136777778888888888888888888888888888888999aab500000100000112238bbbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd153:mariob=956'hfffffffffffffffffffffffffffffffffffffffffc6322343221169998888888887877777777777752011111211112111111111111111112577777778888888888888888888888888888888999aba10000000111011225abacfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd154:mariob=956'hfffffffffffffffffffffffffffffffffffffffffdb96444322110158a998888888887877778885200111111111111111111331111112467777777788888888888888888888888888888888999ab400000000011111248bbaefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd155:mariob=956'hfffffffffffffffffffffffffffffffffffffffffeb99994322211100147899999988888887530011111111111111111111255666677777667777778888888888888888888888888888888899ab800000100011112237ababffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd156:mariob=956'hffffffffffffffffffffffffffffffffffffffffffb9989632221111110011345556665432100111111111111111111111145666677666677777778888888888888888888888888888888889aba20000001111111236abbbdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd157:mariob=956'hffffffffffffffffffffffffffffffffffffffffffda999732221111111111100000000001111111111111111111111111356667776546677777778888888888888888888887887888888899ac50000000111111235abbacfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd158:mariob=956'hffffffffffffffffffffffffffffffffffffffffffeb99895222211111111211111111111111111111111111111111111366677777534567777778888888888888888887877777777888899ab80000011111122347abbabffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd159:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffc99888422211111111221111111111111111111111111111111113666777765356667777778888888888888888877777777777788899ba1010111111222458bbbabfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd160:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffea998872222111111122111111111111111221111111111111114667777764456667777788888888888888888887777777777778889ab301111111223358abbbabefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd161:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffc99988732222111111221111111111111122222221111111136777777644566777777788888888888888888777777777777777888ab30112222334579abbbaacfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd162:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffea9998973222221113532211111111111124432221111123677777764456677777777888888888888888887777777777777777889a523334455678abbbbaabdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd163:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffca99988863211236775222111111111135566666555567777777543566777777777788888888888877887777777777777777789a64567666569bbbbbaabeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd164:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffb9998888887788777763222211111157666677777777777654345677777777777888888888888878777777777777777777778966777532235abbaabceffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd165:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffea999888888887777777632221123556777777777766654445667777777777778888888888887888777777777777777777788556665333347bbbdefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd166:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffca9998888888877777777765567665544555554443344566777778877777778888888888888877777777777777777777787555554433336ababfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd167:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffca999888888888777777777777766666555555666677777888888777777778888888888877777777777777777766677764455443333359bbbdfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd168:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffb99998888888887777777777777777777777777888888888888777777778888888888878777777777777777666667743444443333359bbacffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd169:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffb99988888888888777777777777777788888888888888888777777777888888888878877777777777776666666774444555567778abbbbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd170:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffba9988888888888877777777777788888888888888887777777777788888888888777777777777776666666676445566689aa99aaaabefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd171:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffba99888888888888777777777788888888888888777777666777788888888888877777777777776666666675455566899999999999aefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd172:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffba9998888888888888788787888888888777777777766677788888888888778777777777777766666667644556679999a86545689aadffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd173:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffdaa9998888888888888788888887777777777777666777888888888887787777777777776666666667645566689999520000001257adfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd174:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffeba99888888888888888888887777777777777677778888888888888787777777777777666666677545566799996100000000000136affffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd175:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffcaa999888888888888888888877777777777788888888888888877777777777777766666666764456667999930000000000000001248dfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd176:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffebaa999988888888888888888888888888888888888888888877877777777777666666667654556768999600000000000000000011246aeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd177:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbaa99988888888888888888888888888888888888888888877777777777766666666765566677899a5000000000000000000001112359effffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd178:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbaa9988888888888888888888888888888888888888877777777777776666666765556677789995000000000000000000000001112348dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd179:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbaa9988888888888888888888888888888888888877777777777766666666765566777789994000000000000000000000000001112347cffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd180:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecaa998888888888888888888888888888888788777777777776666666676556667787899a5000000000000000000000000000001112337dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd181:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffca9998888888888888888888888888888777777777777777666666677656667778889996000000000000000000000000000000011112337dffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd182:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeb99988998888888888888888888888887777777777777766666666666566677778889997000000000000000000000000000000000001112348effffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd183:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda9999986589888888888888888888887777777777777776666666666666677778888999810000000000000000000000000000000000001112235afffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd184:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeba99989854434888888888888787777777777777777766666666666665677777888989a9920000000000000000000000000000000000000001112235cfffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd185:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffebaaa99999754431236888887877777777777777777776666666666666666777788888989a9950000000000000000000000000000000000000000001112238efffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd186:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffe968baaa99a755521232027877777777777777777777666666666666666667777788888989a997000000000000000000000000000000000000000000001112235bffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd187:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffc754adbbaaa9655511232100047877777777777766666666666666666666677788888888999aa98100000000000000100100000000000000000000000000000012247effffffffffffffffffffffffffffffffffffffffffffffffff;
10'd188:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffea7544aeccbbba7554112221000001577777777666666666666666666666667777888888999999a9930000000000000000000100000101000000000000000000000012235bfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd189:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffd964443afedccbb8774012221100000002577666666666666666666665566677788888889999999a9970000000000001111110000000100000000000000000000000000112248ffffffffffffffffffffffffffffffffffffffffffffffff;
10'd190:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffb6443332afeeddcb9885012221100000000000356666655555555554456567778888888999999999aa98100000000001111100011011100001000000000000000000000000112235cffffffffffffffffffffffffffffffffffffffffffffff;
10'd191:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffea644333229ffeeedca996112221100000000000000012334443332100366677788888899999999999aa9930000000000111111101000010101000000000000000000000000000011235afffffffffffffffffffffffffffffffffffffffffffff;
10'd192:mariob=956'hffffffffffffffffffffffffffffffffffffffffffff95433222218ffffeeebab61122211000000000000000000000000000003777788888889999999999a9aaaa60000000001111111101110110101010100000000000000000000000000111237ffffffffffffffffffffffffffffffffffffffffffff;
10'd193:mariob=956'hfffffffffffffffffffffffffffffffffffffffffe953322212107ffffffebab70122211100000000000000000000000000004887888888999999999aaaaaabb98000000000001111111110000001101010101001000000000000000000000012225cffffffffffffffffffffffffffffffffffffffffff;
10'd194:mariob=956'hfffffffffffffffffffffffffffffffffffffffea533222111115ffffffebab712222111000000000000000000000000000038888899999999999aaaaaababba940000000000111111110100010101101010101101000000000000000000000011234afffffffffffffffffffffffffffffffffffffffff;
10'd195:mariob=956'hffffffffffffffffffffffffffffffffffffffb6332211111103effffffbbb8112221110000000000000000000000000000199889999999999aaaaaaabbbbcba70000000000001111111100001001111110101010000000000000000000000000011238ffffffffffffffffffffffffffffffffffffffff;
10'd196:mariob=956'hffffffffffffffffffffffffffffffffffffc63322111111102efffffebbb811221111110000000000000000000000000018a999999999aaaaaaaabbbbbbcca9200000000000011111100100001001011111111111110100000000000000000000011236dffffffffffffffffffffffffffffffffffffff;
10'd197:mariob=956'hffffffffffffffffffffffffffffffffffd743222111111100cfffffecbb811222211110000000000000000000000000007baaaaaaaaaaaaaabbbbbccccccba50000000000000111110000000101111011111111111110000000000000000000000101225cfffffffffffffffffffffffffffffffffffff;
10'd198:mariob=956'hfffffffffffffffffffffffffffffffff94322111111111009ffffffbbb911122211111100000000000000000000000004cbbbbbbbbbbbbbbbbccccccccdda91000000000000011110010000000010111111111111111101010100000000000000000111349ffffffffffffffffffffffffffffffffffff;
10'd199:mariob=956'hfffffffffffffffffffffffffffffffa53222111111111008fffffecbb90111221111110100101111000000000000136aedcddddddddddddddddddddddddca500000000000000011110000000010010111111111111110101010100000000000000001111138fffffffffffffffffffffffffffffffffff;
10'd200:mariob=956'hfffffffffffffffffffffffffffffc633221111111111105fffffecbb91011222111111111111111111000001359cefffedeeeeeeeeeeedddddddddddddda81000000000000000110000000000000010111111111111111111010000000000000000000012237efffffffffffffffffffffffffffffffff;
10'd201:mariob=956'hfffffffffffffffffffffffffffe8432211111111111102ffffffcbb800111121111111111110000000147adffffeeeeeeefeb975568aefeeeeeeeeddeeda500000000000000000100000000010001110111111111111111111100100000000000000000111236dffffffffffffffffffffffffffffffff;
10'd202:mariob=956'hffffffffffffffffffffffffffa4322111111111100001cfffffcbbbeda52110000000000012469acefffffffeeeeeeffed844444332236beeeeeeedeeeb81000000000000000000000000000000000010111111111111111111010100000000000000000111125cfffffffffffffffffffffffffffffff;
10'd203:mariob=956'hffffffffffffffffffffffffd73222111111110012342afffffdcbbefffffecba99999abcdeffffffffffffeeeeeeeefe9544333333343347deeeeedeeda600000000000000000000000000000000010111111111111111111111110100000000000000000011224bffffffffffffffffffffffffffffff;
10'd204:mariob=956'hfffffffffffffffffffffffa4222111111110037887779efefdcbbdffffffffffffffffffffffffffffffffffeeeeefe744333333333333445bfeedeeec92000000000000000000000000000000000000011111111111111111111010100000000000000000112234cfffffffffffffffffffffffffffff;
10'd205:mariob=956'hfffffffffffffffffffffd7322111111111027965444448ffeccbdfffffffffffffffffffffffffffffeeeeeeeeeeee64433333333333333344beedeeea700000000000000000000000000000000000000101111111111111111111010101000000000000000011124bffffffffffffffffffffffffffff;
10'd206:mariob=956'hffffffffffffffffffffc43211111111110497543333338feccbcffffffffffffffffffffffffffeeeeeeeeeeeeeef9443333333333333333345dedeeda4000000000000000000000000000000000000000101111111111111111111011101000000000000000111224bfffffffffffffffffffffffffff;
10'd207:mariob=956'hfffffffffffffffffffa32211111111100596443333323cfccbbeeeeeffffffffffffffeeeeeeeeffffffefeeeeefc54333333333333333333337deeec910000000000000000000000000000000000000000101111111111111111111111110000000000000001011235cffffffffffffffffffffffffff;
10'd208:mariob=956'hfffffffffffffffffe6321111111111106954433332328fdccbeffffffffeeeeeeefffffffffffffffffeeeeeeeee843333222223233333333332afeeb6000000000000000000000000000000000000000000110111111111111111111111111000000000000000111225dfffffffffffffffffffffffff;
10'd209:mariob=956'hffffffffffffffffe6321111111111105964433222323deccbeffffffffffffffffffffffffffffffffefeeeeeefc5433325732223333333333425feda40000000000000000000000000000000000000000000000111111111111111111111111000000000000001112237effffffffffffffffffffffff;
10'd210:mariob=956'hfffffffffffffffe5311111111111103964433274231beccbdffffffffffffffffffffffffffffffffefeeeeeeefa433324dfa3233333333333321ced9200000000000000000000000000000000000000000000001011111111111111111111111100000000000000112249ffffffffffffffffffffffff;
10'd211:mariob=956'hffffffffffffffe53111111111111028754322bc3327fdcbcffffffffffffffffffffffffffffffffffeeeeeeeef9433326efa32333333333333309ec9300000000000000000000000000000000000000000000000010111111111111111111111100000000000000101235bfffffffffffffffffffffff;
10'd212:mariob=956'hfffffffffffffe62111111111111006854333494224edcccefffffffffffffffffffffffffffffffffeeeeeeeeee843333367433333333333333308db97000000000000000000000000000000000000000000000000000111111111110111001000000000000000000011237dffffffffffffffffffffff;
10'd213:mariob=956'hfffffffffffff82111111110111103964433332332ceccbeffffffffffffffffffffffffffffffffffffeeeeefee843333322333333333333333308ca9a300000000000000000000000000000000000000000000000000010010000000000000000000000000000000001224aefffffffffffffffffffff;
10'd214:mariob=956'hffffffffffff93110111011011000775433333331bfdccdfffffffffffffffffffffffffffffffffeffeeeeeeeeda43333333333333333333333208ba9b9000000000000000000000000000000000000000000000000000000000000001100000000000000000000000011237bfffffffffffffffffffff;
10'd215:mariob=956'hfffffffffffb31100000000000002865433333317fdccdfffffffffffffffffffffffffffffffffffffeeeeeeeedd4333333333333333333333311ab99cd1000000000000000000000000000000000000000000000000000000000011111000000000000000000000000012259effffffffffffffffffff;
10'd216:mariob=956'hffffffffffd51100000010000000485433333317fdccceffffffffffffffffffffffffffffffffffffefeeeefeede8233333333333333333333204aa99ce6000000000000000000000000000000000000000000000000000000000111111100000000000000000000000011237cffffffffffffffffffff;
10'd217:mariob=956'hffffffffff71101000000000000067543333316eeccceffffffffffffffffffffffffffffffffffffffeeeeffeeeed333333333333333333333018aa99ddc200000000000000000000000000000000000000000000000000000001111111000000000000000000000000000225adfffffffffffffffffff;
10'd218:mariob=956'hfffffffffa3111111100000000017644333314efdccdffffffffffffffffffffffffffffffffffffffeeeeeefeeeee923333233333333333331059ba9adde8000000000000000000000000000000000000000000000000000000111111111000000000000000000000000002238cfffffffffffffffffff;
10'd219:mariob=956'hffffffffe5110111111000000002854333214dfdccdefffffffffffffffffffffffffffffffffffffffeeedbcefeeee7223222222222223321048ac99bdddd400000000000000000000000000000000000000000000000000011111111111000000000000000000000000000236beffffffffffffffffff;
10'd220:mariob=956'hffffffff9210111111100000000285433323dfedccefffffffffffffffffffffffffffffffffffffffeeeeeb9befeeee822222222222222211499bd99bddddc00000000000000000000000000000000000000000000000000111111111111000000000000000000000000000125acffffffffffffffffff;
10'd221:mariob=956'hfffffffe511011111111000000027533322bfedccdffffffffffffffffffffffffffffffffffffffffefeeeec9adfeeeeb312222222222222599bec99cdddde800000000000000000000000000000000000000000000000011111111111110000000000000000000000000000248bffffffffffffffffff;
10'd222:mariob=956'hfffffffa21011111111100000001753322bfecbacffffffffffffffffffffffffffffffffffffffffffeeeeeeea9cefeeeea41112222222589adeea9adddddde70000000000000000000000000000000000000000000000111111111111111000000000000000000000000001228bdfffffffffffffffff;
10'd223:mariob=956'hfffffff62101111111111000000055332afeba9beffffffffffffffffffffffffffffffffffffffefffeeeeeeeeb9befeeeeec8543345789aceeeea9addcddddd5000000000000000000000000000000000000000000001111111111111110000000000000000000000000000136acfffffffffffffffff;
10'd224:mariob=956'hffffffc41101111111111100000036429feba9bfffffffffffffffffffffffffffffffffffffffffffeefeeeeeeec9adeeeedeeeeddddddeeeeeee99bddddddddd300000000000000000000000000000000000000000011111111111111111000000000000000000000000000125abfffffffffffffffff;
10'd225:mariob=956'hffffff9310011111111111100000076bfdb99dfffffffffffffffffffffffffffffffffffffffffffeffeeeeeeeeeea9ceeeeeeeeeefffeeeeeddc99ceddcdddddd40000000000000000000000000000000000000000111111111111111111000000000000000000000000000025abeffffffffffffffff;
10'd226:mariob=956'hffffff62100111111111111100008eefdbaaeffffffffffffffffffffffffffffffffeffffffffffeeefeefeeeeeeeeb9bdeeeeeeeddccbbaaaaaa9acddddcdddddd40000000000000000000000000000000000000011111111111111111111000000000000000000000000001249beffffffffffffffff;
10'd227:mariob=956'hfffffe5110011111111111111104effdb99efffffffffffffffffffffffffffffffffffffeffffefeefeefeeeeeeeeeed9acccbbaaaa9a999998889addddddcdddddd300000000000000000000000000000000000011111111111111111111110000000000000000000000001125aadffffffffffffffff;
10'd228:mariob=956'hfffffd3100011111111111111106ffdb9aeffffffffffffffffffffffffffffffeffffffffeffefeefefeeeeeeeeeeeeeea9999998888888888999abeddddddcddddde60000000000000000000000000011000000111111111111111111111111000000000000000000000000125aadffffffffffffffff;
10'd229:mariob=956'hfffffb2100011111111111111105febaaeffffffffffffffffffffffffffffffffffffffffffefffeefeefeeeeeeeeeeeeec988999aabccdddddddddddddddddcdddddd9000000000000000000000000133200001111111111111111111111110000000000000000000000001126aadffffffffffffffff;
10'd230:mariob=956'hfffffa2100001111111111111104ecaaeffffffffffffffffffffffffffffffffeffffffefeeeefeeeeeeeeeeeeeeeeeeeeedccdeeeeeeeeeeeeeeeedddddddddcdddddeb10000000000000000000002443000011111111111111111111111101000000000000000000000000137badffffffffffffffff;
10'd231:mariob=956'hfffff921000011111111111111117aaeffffffffffeffeefefffffffffffffffffeffeeefeffffeeeefeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddcddddddd7000000000000000000155530000111111111111111111111110000000000000000000000000001238baeffffffffffffffff;
10'd232:mariob=956'hfffff821000011111111111111104bdffffeffeffffeefffeefffeffeffffffefeffefefefeefeefefeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddccdddddcdb40000000000000005ab8400001111111111111111111111110000000000000000000000000001249bbeffffffffffffffff;
10'd233:mariob=956'hfffff82100001111111111111111afffffeefffefeffeeeeefefefefefffefefefeefefeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddccdddcccdda40000000000058bc9610000111111111111111111111101000000000000000000000000001226abbfffffffffffffffff;
10'd234:mariob=956'hfffff82100000111111111111104effffeeefeeffeefffefeeeefefffefeffffeffeefeeeefeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddcdddcccccdd952111257adc787100011111111111111111111111100000000000000000000000000001238bbcfffffffffffffffff;
10'd235:mariob=956'hfffff8210000001111111111110affffeefeeefeeefeeeeeefffefffefefeffefefeeeefefeeeefeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddccdccccccccccbbbbbb89999300001111111111111111111111100000000000000000000000000001125abadfffffffffffffffff;
10'd236:mariob=956'hfffff8210000011111111111112effefefeefeeeeeeefeeeeefefeffeffffeefefeefefefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdddddddddddddcccccccccbbbbbaaa989996000011111111111111111111111100000000000000000000000000001236bbbefffffffffffffffff;
10'd237:mariob=956'hfffff8210000001111111111107fefeeefeeeeeeeeeeeefefefeeeeefeeeeefefeefeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeededddddddddddddcdcccccccccbbbbbaaa99a881000111111111111111111111110000000000000000000000000000011259bacffffffffffffffffff;
10'd238:mariob=956'hfffff921000001111111111111cffeeeeeeeeeeeeeeeeeeeefefeeefeeefeeeefeeeeeeeefeeeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddcdcccbccccbbbbbaaa99984000111111111111111111111110000000000000000000000000000001237abbdffffffffffffffffff;
10'd239:mariob=956'hfffffa21100000111111111114efeeeeeeeeeeeeeeeeeeeeeeeeeefeeefeeeefeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeededdeddddddddddddcdccccccbbbbbbbaaa99aa70001111111111111111111111100000000000000000000000000000012249bbbfffffffffffffffffff;
10'd240:mariob=956'hfffffb31000000011111111118ffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddcdccccccccbbbbaaaaa99992000111111111111111111111100000000000000000000000000000001237bbadfffffffffffffffffff;
10'd241:mariob=956'hfffffd3110000001111111111bfeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddddccccccccccbbbbaaa999a6000111111111111111111111100000000000000000000000000000001225abbbffffffffffffffffffff;
10'd242:mariob=956'hfffffe5210000000111111113efeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdededdddddddddddcdccccccccbbbbaaabbbba2001111111111111111111110000000000000000000000000000000001248bbadffffffffffffffffffff;
10'd243:mariob=956'hffffff6210000000111111107feeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdedddddddddddddddddcccccccbbbbabddddde7000111111111111111111110000000000000000000000000000000001236abacfffffffffffffffffffff;
10'd244:mariob=956'hffffff821100000011111110afeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdedddddddddddddddddccccccccbbbaceeddddb100111111111111111111111000000000000000000000000000000001235abbbefffffffffffffffffffff;
10'd245:mariob=956'hffffffa31000000001111111cfeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededeededddddddddddddddcdccccbcbbbaceeeeedd5001111111111111111111111000000000000000000000000000000001248bbadffffffffffffffffffffff;
10'd246:mariob=956'hffffffc42100000000111113efeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeededddddddddddddddddcdccccccbbbbceeeeeeea110111111111111111111110100000000000000000000000000000001237bbabfffffffffffffffffffffff;
10'd247:mariob=956'hffffffe62100000000111105feeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddddddcdccccccbbbbbeeffeeee910111111111111111111111000000000000000000000000000000001236abbbefffffffffffffffffffffff;
10'd248:mariob=956'hfffffff92110000000111108feeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddddddcdcdccccbbbbacefffffee90011111111111111111111100000000000000000000000000000001134abbadffffffffffffffffffffffff;
10'd249:mariob=956'hfffffffb421000000001100afeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdeddddddddddddddccccccbbbbaaeffffffffb1011111111111111111111000000000000000000000000000000012349bbacfffffffffffffffffffffffff;
10'd250:mariob=956'hfffffffe521000000000018eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdeddddddddddddddcdccccccbbbabeffffffffe401111111111111111111000000000000000000000000000000012248bbabffffffffffffffffffffffffff;
10'd251:mariob=956'hffffffff8221000000005ffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededededddddddddddddddcdccccccbbbaabffffffffffa0111111111111111111000000000000000000000000000000012247bbabeffffffffffffffffffffffffff;
10'd252:mariob=956'hffffffffc3210000002bfffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdeddddddddddddddcdcccccccbbbbacfffffffffff601111111111111111100000000000000000000000000000011237bbbbefffffffffffffffffffffffffff;
10'd253:mariob=956'hfffffffff621000004effffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdeddddddddddddddcdcdcccccbbbbaabfffffffffffe4011111111111111110000000000000000000000000000011236abbadffffffffffffffffffffffffffff;
10'd254:mariob=956'hfffffffff93210007ffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddddddddddccccccccbbbbaabefffffffffffe40111111111111111000000000000000000000000000111236abbadfffffffffffffffffffffffffffff;
10'd255:mariob=956'hfffffffffc42100bffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdeddddddddddddddddcdcccccccbbaa998effffffffffffe301111111111111100000000000000000000000000111236abbacffffffffffffffffffffffffffffff;
10'd256:mariob=956'hffffffffff7211bfffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdededdddddddddddddddcdcccbbaa99999adfffffffffffffe4011111111111100000000000000000000000000012236abbacfffffffffffffffffffffffffffffff;
10'd257:mariob=956'hffffffffffa32cfffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededeededddddddddddddcccbbaaaabbbbcccccaceffffffffffffff60111111111110000000000000000000000000012336abbacffffffffffffffffffffffffffffffff;
10'd258:mariob=956'hffffffffffd5cffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdededddddddccbbbbbbbcccdddddcccbbbbaaceeffffffffffffff811111111110100000000000000000000000112336abbacfffffffffffffffffffffffffffffffff;
10'd259:mariob=956'hfffffffffffdffffffeeedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddcccbbbbbccdddddeddddddcccccbbbbaaaedefffffffffffffffa101111111000000000000000000000000012336abbacffffffffffffffffffffffffffffffffff;
10'd260:mariob=956'hffffffffffffffffeeeddcdeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddccccbbbbcccddeeeeeeeeddddddddcccccccbbbbaa9cfedefffffffffffffffe3011101000000000000000000000000012336abbacfffffffffffffffffffffffffffffffffff;
10'd261:mariob=956'hfffffffffffffffeeeddcdeccdeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddcccbcbcccddddeeeeeeeeeeedddddddddddcdcccccccbbbbababeefddeffffffffffffffff70011000000000000000000000000112346abbacffffffffffffffffffffffffffffffffffff;
10'd262:mariob=956'hffffffffffffffeeeddcbdffdcbbccddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddcccbbbbbcccdddeeeeeeffeeeeeeeeededdddddddddddddcdcccccccbcbbbbaabffefddeefffffffffffffffc10000000000000000000000000012246abbacfffffffffffffffffffffffffffffffffffff;
10'd263:mariob=956'hfffffffffffffeeedccbadeefffeedccbbbbbbccccccccccccccccccccccccbcbbbbbbbbcccdddeeeffffffffeeeeeeeeeeeedeededdddddddddddddddcdcdcccccbcbbbbaaadeffffcceeffffffffffffffff700000000000000000000000012247abbacffffffffffffffffffffffffffffffffffffff;
10'd264:mariob=956'hfffffffffffeeeedccbbdeeeeeeefffffeeeeeddddddddddddddddddddeeeeeeeeeeeffffffffefeeeeeeeeeeeeeeeeeeeeedddddddddddddddddddddddcdcccccccbbbbbb9cefefffecceeefffffffffffffffc300000000000000000000012247abbacfffffffffffffffffffffffffffffffffffffff;
10'd265:mariob=956'hffffffffffeeeedcbbbdfeeeeeeeeeeeeeeeeeffffffffffffffffffffffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddddddddcdcdcccccccbcbbbbaaceeffffffccdeeefffffffffffffff9100000000000000000011247abbacffffffffffffffffffffffffffffffffffffffff;
10'd266:mariob=956'hfffffffffeeeddcbbbdffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeeeedededddddddddddddddddddddcdcdcdcccccbbbbbbaa9efffffffffccdeeeeeffffffffffffff9100000000000000001238bbbacfffffffffffffffffffffffffffffffffffffffff;
10'd267:mariob=956'hfffffffffeeedcbbbcfffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeededededddddddddddddddddddcdcdcdcccccbbbbaaaa9aeefffffffffccdeeeeeeeefffffffffffe9200000000000001236cbbacffffffffffffffffffffffffffffffffffffffffff;
10'd268:mariob=956'hfffffffffeedccbbbffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeeeeeedededeededddedddddddddddddddddddcdcdccccbbbbaaaaa9999befffffffffffcbcdeeeeeeeeeeffffffffffb4000000000011249bcbdfffffffffffffffffffffffffffffffffffffffffff;
10'd269:mariob=956'hfffffffffedccbbbfffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeeeeeedeeeeeedededeedededdddddddddddddddcdcccccccbbbbabbbbccdcabbaadeffffffffffffdbcddeeeeeeeeeeeefffffffffa400000001148acdbefffffffffffffffffffffffffffffffffffffffffff;
10'd270:mariob=956'hfffffffffedcbbbefffffeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeeeeeeeeeedeeeeeededeeeededeeeddeddddddddddddddddccccbbbbbbbcccdddddddccbaabaaaeefffffffffffffdbccddeeeeeeeeeeeeeffffffffeb84322369abcccbfffffffffffffffffffffffffffffffffffffffffff;
10'd271:mariob=956'hfffffffffeccbbcffffffeddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededeeeeeedededeedededdddddddddddddccccbbbbbbccddddededddddccccbcbbabab9beeffffffffffffffebbccdddeeeeeeeeeeeeeffffffffffffffeedccdbdffffffffffffffffffffffffffffffffffffffffff;
10'd272:mariob=956'hfffffffffecbbbffffffffdcddddeddeeeeeeeeeeeeeeeeeeedededededeeeededededdddededdddddddddddddccccbcbcccccdddeeeeeeeddddcdcccccccccccbbaabbaabefffffffffffffffffcbbccddddddddeddeeeeeeeeffffffffeeeeeedbbffffffffffffffffffffffffffffffffffffffffff;
10'd273:mariob=956'hffffffffffdcbefffffffeeedcccdddddddddddddedddeddddededddddddddddddddddddddddddddcdccccccccccdddeeeeeeeeedddddddcdddcdcccccccccccbbbaabaa9ceefffffffffffffffffcbbcccdddddddddddddeeeeeeeeeeeeeeeeeedbbefffffffffffffffffffffffffffffffffffffffff;
10'd274:mariob=956'hfffffffffffcdffffffffeeeffedccccccccdddddddddddddddddddddddddddddcccccccccbcbcccccdddeeeeeeeeeeeddddddddddddddcdcdcdccccccccccccbbbaabaaadefffffffffffffffffffeaabccccdddddddddddddddeeeeeeeeeeedddbaefffffffffffffffffffffffffffffffffffffffff;
10'd275:mariob=956'hffffffffffffffffffffffeeedeefffeedddccccccccccccccccccbcbcbccccccccdddedeeeeffffeeeeeeeddddddddddddddddddddddddddccccccccccccccbbbbaaaaaadeeffffffffffffffffffffc9abbccccccccccccccddddddddddddccdcabefffffffffffffffffffffffffffffffffffffffff;
10'd276:mariob=956'hffffffffffffffffffffffeeeeedeeeeeeeeeffeeeeeeeeeeeeeeeeeeefeefffffeeeeeeeeeeddeddddddddddddddddddddddddddddddcdddcccccccccccccbbbbbaaaaaadeffffffffffffffffffffffeb9abbbbccccccccccccccccccccccccdbbbefffffffffffffffffffffffffffffffffffffffff;
10'd277:mariob=956'hffffffffffffffffffffffeeeededddddddddddeeeeeeeeeeeeeeedeeeeddddddddddddddddddddddddeddddddddddddddddddddddcdddcccdcccccccccccbbbbbbaaaa9aeeffffffffffffffffffffffffda9abbbbbbbccccccccccccccccccdcbbbffffffffffffffffffffffffffffffffffffffffff;
10'd278:mariob=956'hffffffffffffffffffffffedeeeedddddddddddddddddddddddddddddddddddddededddedddddddddddddddddddddddddddddddddcdcdcdcdccccccccccccbbbbbbaaaa9beefffffffffffffffffffffffffeba99abbbbbbbbcccccccccccccccbbacffffffffffffffffffffffffffffffffffffffffff;
10'd279:mariob=956'hffffffffffffffffffffffedededdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcccccccccccccccccccbbbbbbaaaaa9beefffffffffffffffffffffffffeeca989abbbbbbbccccccccccccdbbbbeffffffffffffffffffffffffffffffffffffffffff;
10'd280:mariob=956'hffffffffffffffffffffffedddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddccccccccccccccccccbcbbbbbbbaaaa9beefffffffffffffffffffffffffeeecaa889aabbbbbbbccccccccddcaadfffffffffffffffffffffffffffffffffffffffffff;
10'd281:mariob=956'hffffffffffffffffffffffeddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddccccccccccccccccccbbbbbbbbbaa9999ceefffffffffffffffffffffffffeeedcaaaa999aaabbbbbbbccccdddbcffffffffffffffffffffffffffffffffffffffffffff;
10'd282:mariob=956'hfffffffffffffffffffffffddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddccccccccccccccccccccbbbbbbbbaaa9998ceefffffffffffffffffffffffffeeeddbbaaaaaaaaaaaabbbbcccdddbcffffffffffffffffffffffffffffffffffffffffffff;
10'd283:mariob=956'hfffffffffffffffffffffffdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcccccccccccccccccccbbbbbbbbbbaaaa998ceefffffffffffffffffffffffffeeeddcbbbbaaaaaaabbbbbccccdddbbffffffffffffffffffffffffffffffffffffffffffff;
10'd284:mariob=956'hfffffffffffffffffffffffedddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcccccccccccccccccccccbbbbbbbbbbaaaaa998ceefffffffffffffffffffffffffeeeddcbbbbbbbbbbbbbbbcccccddecaefffffffffffffffffffffffffffffffffffffffffff;
10'd285:mariob=956'hfffffffffffffffffffffffeddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcccccccccccccccccccbcbbbbbbbbbbbaaaaa998ceefffffffffffffffffffffffffeeeddcccbbbbbbbbbbbbbccccccddcadfffffffffffffffffffffffffffffffffffffffffff;
10'd286:mariob=956'hfffffffffffffffffffffffeddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddccccccccccccccccccccccbbbbbbbbbbabaaaa9998ceeefffffffffffffffffffffffeeeeddcccbbbbbbbbbbbbcccccccdddbcfffffffffffffffffffffffffffffffffffffffffff;
10'd287:mariob=956'hffffffffffffffffffffffffddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddccccccccccccccccccccbbbbbbbbbbbbbbbbaaaa9988ceeefffffffffffffffffffffffeeeeddccccbbbbbbbbbbbcccccccdddbbfffffffffffffffffffffffffffffffffffffffffff;
10'd288:mariob=956'hffffffffffffffffffffffefedddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddccccccccccccccccccccccbbcbbbbbbbbbbbbaaaaaa99988ceeefffffffffffffffffffffffeeeeddcccccbbbbbbbbbbcccccccdddbbfffffffffffffffffffffffffffffffffffffffffff;
10'd289:mariob=956'hfffffffffffffffffffffefeeddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddcdccccccccccccccccbcccbbbbbbbbbbbbbbbbaaaaa998887ceeeffffffffffffffffffffffeeeeeddccccccbbbbbbbbbbccccccdddcbeffffffffffffffffffffffffffffffffffffffffff;
10'd290:mariob=956'hffffffffffffffffffffffeeeddddddddddddddddddddddddddddddcdddddcddddddddddddddddddddddcdccccccccccccccccccbcbbbbbbbbbbbbbbbbbbaaaaa999a9aaceeefffffffffffffffffffffeeeeedddcccccccbbbbbbbbbcccccccdddadffffffffffffffffffffffffffffffffffffffffff;
10'd291:mariob=956'hfffffffffffffffffffffeeeeeddddddddddddddddddddcddcddcdddcdcdddcdcdddddddddddddddddccdccccccccccccccccccbbbbbbbbbbbbbbbbbbbbaaaaaaabcccccdeeefffffffffffffffffffffeeeeeddcccccccccbbbbbbbbbbccccccddbcffffffffffffffffffffffffffffffffffffffffff;
10'd292:mariob=956'hfffffffffffffffffffffeeeeedddcdcddcdddccddddcdcddddcdcccccdcdcdcdcdccdddcdddccdcdcccccccccccccccccccbbbbbbbbbbbbbbbbbbbbbbbbbbbccdddddccdeeeefffffffffffffffffffeeeeeeddccccccccbbbbbbbbbbbbcccccddbbffffffffffffffffffffffffffffffffffffffffff;
10'd293:mariob=956'hffffffffffffffffffffeeeeeeeddcccccdccddccdccccccdccdcccccdccccccccccdccccccccccccccccccccccccccccbbbbbbbbbbbbbbbbbbbbbbbbbbcccdddddddddcdeeeefffffffffffffffffffeeeeeeddccccccccbbbbbbbbbbbbccccccdcbefffffffffffffffffffffffffffffffffffffffff;
10'd294:mariob=956'hfffffffffffffffffffffeeeeeedcccccccccccccccccdcccccccccccccccccccccccccccccccccccccccccccccccccccbbbbbbbbbbbbbbbbbbbbbbbbbcccdddddddddccdeeeeffffffffffffffffffeeeeeedddcccccccccbbbbbbbbbbbccccccddbdfffffffffffffffffffffffffffffffffffffffff;
10'd295:mariob=956'hffffffffffffffffffffeeeeeeedccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccbbbbbbbbbbbbbbbbbbbbbcbbccccdddddddddddddcceeeeffffffffffffffffffeeeeeeddccccccccccbbbbbbbbbbbcccccccdbbfffffffffffffffffffffffffffffffffffffffff;
10'd296:mariob=956'hfffffffffffffffffffffeeeeeeedccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccbbbbbbbbbbbbbbbbbbbbbbbcccccddddddddddddddcddeeeffffffffffffffffeeeeeeeeddccccccccccbbbbaabbbbbcccccccdcbfffffffffffffffffffffffffffffffffffffffff;
10'd297:mariob=956'hffffffffffffffffffffeeeeeeeedccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccbbbbbbbbbbbbbbbbbbcbbccccdddddddeddddddddcdcdeeefffffffffffffffffeeeeeedddccccccccccbbbaaaabbbbbcbcccccdbdffffffffffffffffffffffffffffffffffffffff;
10'd298:mariob=956'hfffffffffffffffffffefeeeeeeeeccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccbbbbbbbbbbbbbbbbbbbbbbcccddddddddeddeddddddddcdeeefffffffffffffffeeeeeeeeddcccccccccccbbaaaaabbbbbbbbccccddbffffffffffffffffffffffffffffffffffffffff;
10'd299:mariob=956'hfffffffffffffffffffeeeeeeeeeedcccccccccccccccccccccccccccccccccccccccccccccccccccccccccccbbbbbbbbbbbbbbbbbbbbbbcccdddddddddeededdddddddccdeeeeffffffffffffffeeeeeeedddcccccccccccbbaaaaabbbbbbbbbcccddbdfffffffffffffffffffffffffffffffffffffff;
10'd300:mariob=956'hfffffffffffffffffffffeeeeeeeeecccccccccccccccccccccccccccccccccccccccccccccccccccccccccccbbbbbbbbbbbbbbbbbbbbccccddddddedeeededdedddddddcceeeeeffffffffffffeeeeeeedddcccccccccccbbbbaaaaaaaabbbbbbcccddcfffffffffffffffffffffffffffffffffffffff;
10'd301:mariob=956'hfffffffffffefffffffeeeeeeeeeeedccccccccccccccccccbcbbbbbbbbcccccbcccccccccccccccccccbccbbbbbbbbbbbbbbbbbbbbccccddddeddeeeeeeeededdddddddcddeeeeffffffffffffeeeeeeedddcccccccccccbbbbaaaaaaaaaabbbbccccdcdffffffffffffffffffffffffffffffffffffff;
10'd302:mariob=956'hfffffffffffeffffffffeeeeeeeeeedcbbcbcbccccccccccbccccccccccccbbbcbcccccccccccccccccbcbbbbbbbbbbbbbbbbbbbbcccccddddddeeeeeeeeededdddddddcdcdeeeefffffffffffeeeeeeeeddcccccccccccbbbbaaaaaaaaaaaabbbbcccddbffffffffffffffffffffffffffffffffffffff;
10'd303:mariob=956'hfffffffffffefffffffeeeeeeeeeeeddbbbbbbbbcbbbbbbbcbbcbbbbbbbbcbbbbcbbbbcbcbccbcbcbccbbbbbbbbbbbbbbbbbbbbbccccdddddddeeeeeeeeedeededddddddccdeeeeeffffffffffeeeeeeeddccccccccccccbbbbaaaaaaa9aaaabbbbccccdcdfffffffffffffffffffffffffffffffffffff;
10'd304:mariob=956'hfffffffffffeefffffefeeeeeeeeeeddcbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbcbcbbbbbbbbbbbbbbbbbbbbaaaaabbbbcccdddddeddeeeeeeeeeeeededdddddddccdeeeeeefffffffeeeeeeeeddcccccccccccbbbbbbacca99999aaaabbbccccddceffffffffffffffffffffffffffffffffffff;
10'd305:mariob=956'hfffffffffffeeeeffffeeeeeeeeeeedddcbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbabaaaaaaabbbbbcdddddeedeeeeeeeeeeeeeeddedddddddcceeeeeffffffffeeeeeeedddccccccccccbbbbbbbbbba999999aaabbbbccccdddffffffffffffffffffffffffffffffffffff;
10'd306:mariob=956'hffffffffffffeeffffeeeeeeeeeeeedddcbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbaaaaaaaaaabbbcccdddddeddeeeeeeeeeeeeeeededddddddcccdeeeefefffffeeeeeeedddccccccccbcbbbbbbbbbbb98889999aaabbbbccccdcefffffffffffffffffffffffffffffffffff;
10'd307:mariob=956'hffffffffffffeeeeeffeeeeeeeeeeedddccbbbaaaaababbababbabababaababbbbbbbbbbbbbbbbbbbbbbaaaaaaaaaaaaaabbcccdddddedeeeeeeeeeeeeeeeededdddddddddcdeeeeeeeffeeeeeeeedddccccccccbbbbbaababbbacb9aa9999aaaabbbcccccdcfffffffffffffffffffffffffffffffffff;
10'd308:mariob=956'hfffffffffffeeeeeffeeeeeeeeeeeedddccbbbbaaaaaaaaaaaaaaabaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbccdddddeeeeeeeeeeeeeeeeeeeeeededddddddccddeeeeeffefeeeeeedddcccccccccbbbbaaaaaababefffffec99aabbbbcccccdddffffffffffffffffffffffffffffffffff;
10'd309:mariob=956'hffffffffffeeddeeefefeeeeeeeeeedddcccbaabbaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabccdddddeeddeeeeeeeeeeeeeeeeeededddddddddccdeeeeeeeeeeeeeedddcccccccccbbbbaaaaaaaacfffffffffdaabbcbbbcccccdcdfffffffffffffffffffffffffffffffff;
10'd310:mariob=956'hffffffffffeedceeeeeeeeeeeeeeeddddcccbaaaabaaaaaaaaaaaaabaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabccdddddeeddeeeeeeeeeeeeeeeeeededeedddddddccdeeeeeeeeeeeeedddccccccccbbbaaa9999aaaafffffffffffdabbbccbbcccccdbfffffffffffffffffffffffffffffffff;
10'd311:mariob=956'hfffffffffeedefeeeeeeeeeeeeeeeddddccccbbaaaaaaaaaaaaaaaaabaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabccdddddddeeeeeeeeeeeeeeeeeeeeeeeeedddddddcccdeeeeeeeeeeeedddccccccccbbbba9988889a9dffffffffffeebbbccccbbccccdccffffffffffffffffffffffffffffffff;
10'd312:mariob=956'hffffffffeeeffffeeeeeeeeeeeeeeddddccbccbaaaabaaaaaaaaaaaaabaaaaaaabaaaaaaaaaaaaaaaaaaaaaaaaaaaaaccdddddeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddddccdeeeeeeeeeeddddcccccccbbbaa988777898aeffffffffffedcddddddbbccccdcbefffffffffffffffffffffffffffffff;
10'd313:mariob=956'hffffffffffffffffeeeeeeeeeeeeedddcccbcccbaaaaaaaaaaaaaaaaaabaaaaaaabaaaaaaaaaaaaaaaaaaaaaaaaaaabcdddddddeeeeeeeeeeeeeeeeeeeeeeeeeededddddddcccdeeeeeeeeeddddccccccbbbbaa9877677788cffffffffffedcdeeeeedcbbbccccadfffffffffffffffffffffffffffffff;
10'd314:mariob=956'hfffffffffffffffffeeeeeeeeeeeddddccbbbdcbaabaaaaaaaaaaaaaaaaaaaaaaaabaaaaaaaaaaaaaaaaaaaaaaaaabcddddddeedeeeeeeeeeeeeeeeeeeeeeeeeeedddddddddcccdeeeeeeeedddccccccbbbaa998766666779efffffffffeedcdfeeedccbbbccccbbfffffffffffffffffffffffffffffff;
10'd315:mariob=956'hffffffffffffffffffeeeeeeeeeddddccbbaacdcbbaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabccddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeddedddddddcccdeeeeeeedddccccbbbbb98887765666678afffffffffeedccceeedccbbbbbcccabeffffffffffffffffffffffffffffff;
10'd316:mariob=956'hfffffffffffffffffffffeeeeeedddccbbaa9cddcbaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabcdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddccccdeeeeedddccbbbcccccb7667775445678cfffffffeeedcccabdcbccbbbbbccbbbeffffffffffffffffffffffffffffff;
10'd317:mariob=956'hfffffeeffffffffffffffeeeeedddccbbaa99bdddcbaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa99a99aaaaaaaabcdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddcccbdeeeeedddccccccccccca889998657779effffffeeeddcccabbbccbaabbccbbbbfffffffffffffffffffffffffffffff;
10'd318:mariob=956'hffffffeeefffffffffffeeeeeeddccbbaaa98addddbbaaaaaaaaaaaa999aaaaaaaaaaaaaaaaa99999999aaaaaaabccddddddeddeeeeeeeeeeeeeeeeeeeeeeeeeedeeddddddddcccbdeeeeeedeeeeeeeedccb99999888888aefffffeeeddcccbabbbccbbbbbbbbbadfffffffffffffffffffffffffffffff;
10'd319:mariob=956'hffffffedeeefffffffffeeeeeddccbbaaa9989ddddcbbaaaaaaaaaaaa99999aaa9aa9aa99a999999999999aaaaabcdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddddcccbceeeeeeeeeeeeeeeeeca88999889999cffffeeeeedccccbbbbbcbbbbbbbbaacffffffffffffffffffffffffffffffff;
10'd320:mariob=956'hfffffffddeeeeeeeeeeeeeeeddcbbaaaaa9989dddddcbbaaaaaaaaaaaa9999889999a999999999999999899aaaabcdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddcccbdeeeeeeeeffffeeedeedb99889999beeffeeeedddcccbabbbccbbbaaaabcefffffffffffffffffffffffffffffffff;
10'd321:mariob=956'hffffffffcddeeeeeeeedddddcbbbaaaaa99989ddddddcbaaaaaaaaaaaaaa999877889999999999999998889aaaabcdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeededdeddddddccccbcdeeeeeeffffffeefffffec87899aefeeeeeeeddccccbbbbccbbabccdeffffffffffffffffffffffffffffffffffff;
10'd322:mariob=956'hffffffffeccdddddddddccbbbbbaaaaaa99aaacddddddcbbaaaaaaaaaaaaaa9998888889999999999988899aaaabccdddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddcccbcdeeeeeeffffffffffffffdceffffffeeeeeddccccbbbbbcbbbbeffffffffffffffffffffffffffffffffffffffff;
10'd323:mariob=956'hfffffffffecccccdcccbbbbbbbbaaaaaaaaaaacdddddddcbbaaaaaaaaaaaaaa9999998888888888888888899aaabcdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddccccbbddeeeeeffffffffffffffffffffffffeedddcccccbbbbcbbbbdfffffffffffffffffffffffffffffffffffffffff;
10'd324:mariob=956'hffffffffffebcccbbbbbbbbbbbbbbbbbaaaaaacddddddddccbaaaaaaaaaaaaaaa9999999988888878888889aaaacccddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddcccccabdeeeeefffffffffffffffffffffffffdddccbccbbbbccaabcefffffffffffffffffffffffffffffffffffffffff;
10'd325:mariob=956'hffffffffffffcbbcbbbbbbbbbbbcbbaaaaaabbcddddddddddcbaaaaaaaaaaaaaaa9999999998888877776669aaabdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddccccc9cddeeeeefffffffffffffffffffffffeccbbbccbbbbcaaabbceffffffffffffffffffffffffffffffffffffffff;
10'd326:mariob=956'hfffffffffffffdbbbbbbbbbbbbbbbbbbbbbbbbbdddddddddddcbbaaaaaaaaaaaaa9999999998888887777667aaabdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddddddccccb8cddeeeefffffffffffffffffffffffedbbbbcbbbbbbaaabbbcefffffffffffffffffffffffffffffffffffffff;
10'd327:mariob=956'hfffffffffffffffdbaaabbbbbaaaaabbbbbbbabddddddddddddccbaaaaaaaaaaaaa9999999998888887777668aacccdddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddccccc98cddeeeeeffffffffffffffffffffeeebbbcbabbbb9aaabbbbcdffffffffffffffffffffffffffffffffffffff;
10'd328:mariob=956'hfffffffffffffffffecbbaabbbcdeecbaaaabbceddddddddddddccbaaaaaaaaaaaaa9999999998888887777669abcddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddccccb79cdddeeeeefffffffffffffffffeeeecbcbabbba9aaabbbbbccdfffffffffffffffffffffffffffffffffffff;
10'd329:mariob=956'hfffffffffffffffffffffeeeffffffffeeeefffeddddddddddddddcbaaaaaaaaaaaa99999999988888877776679bccddddddddddeedeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddddcccca69ccdddeeeeefffffffffffffeeeeedcbbabba99aaabbbbbccccdffffffffffffffffffffffffffffffffffff;
10'd330:mariob=956'hfffffffffffffffffffffffffffffffffffffffedddddddddddddddcbbaaaaaaaaaaa9999999998888887777667bccddddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddccccc878bccdddeeeeefffffffeeeeeeeddccaaba9999aaaabbbbccccbefffffffffffffffffffffffffffffffffff;
10'd331:mariob=956'hfffffffffffffffffffffffffffffffffffffffeddddddddddddddddccbaaaaaaaaaaa9999999988888877777669cccdddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddddddccccb778abccdddeeeeeeeeeeeeeedddccccba98999aaaaabbbccccdbbfffffffffffffffffffffffffffffffffff;
10'd332:mariob=956'hfffffffffffffffffffffffffffffffffffffffeddddddddddddddddddcbbaaaaaaaa99999999998888887777766bccdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddccccc97779bbccdddeeeeeeeeddddcccccc988899999aaabbbbbcccccaeffffffffffffffffffffffffffffffffff;
10'd333:mariob=956'hffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddccbaaaaaaaa99999999988888877777768cccddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddccccb88777abbcccddddddddccccbbbbc988999999aaaaabbbbcccccadffffffffffffffffffffffffffffffffff;
10'd334:mariob=956'hffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddccbaaaaaaa999999999888888777777769ccdddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddddcccca888778abbbbccccccbbbbbbbcb98888999999aaaabbbbcccccacffffffffffffffffffffffffffffffffff;
10'd335:mariob=956'hffffffffffffffffffffffffffffffffffffffffdddddddddddddddddddddccbaaaaaaa99999999888888877777767bcddddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddcdccc98888888abbbbbbbbbbbbbbbbaaaa999999999aaabbbbbcccbacffffffffffffffffffffffffffffffffff;
10'd336:mariob=956'hffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddcbbaaaa9999999998888888777777768ccdddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddccccb9888888889aabbbbbbbbbbbbbaabbaa9999999aaabbbbcccbacffffffffffffffffffffffffffffffffff;
10'd337:mariob=956'hffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddccbbaaaa999999999888888877777777bccdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddcccca8888888888888abbbbbbbaabcdcbbaaaa9999aaaabbbbcbbacffffffffffffffffffffffffffffffffff;
10'd338:mariob=956'hffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddcccbaa99999999998888888777777779ccdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddcdccca9999898999889bbaaaabcdfffffedbaaaaaaaaaabbbbbbbadffffffffffffffffffffffffffffffffff;
10'd339:mariob=956'hffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddcccbaa9999999998888888877777778acdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddccccc9999999999999bbceeffffffffffffedbaabbbbbbbbbbbabfffffffffffffffffffffffffffffffffff;
10'd340:mariob=956'hfffffffffffffffffffffffffffffffffffffffffddddddddddddddddddddddddcdccbaa9999999988888888777777787ccdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddcccb999999999999abcfffffffffffffffffecbbaabbbbbaacffffffffffffffffffffffffffffffffffff;
10'd341:mariob=956'hfffffffffffffffffffffffffffffffffffffffffdddddddddddddddddddddddcdccccbaa999999988888888777777787accdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddcdccca99999999999abbffffffffffffffffffffedcbbbbbcefffffffffffffffffffffffffffffffffffff;
10'd342:mariob=956'hfffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddcdccccbba999999988888887777777878cddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeededeeddddddddddddcdca9999999999abbdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd343:mariob=956'hfffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddcdccccbba99999988888887777777877acddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddcccc999999999aabacffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd344:mariob=956'hfffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddcdcdccccbba99999988888888777778878ccdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddddddcdcb99a99999aaabbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd345:mariob=956'hfffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddccccccbba9999988888888877778877acddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddcccbaaaaa9aaaabbefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd346:mariob=956'hfffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddccccccccbba9999888888888877788778cdddddddddededeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddccccaaaaaaaaaabbcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd347:mariob=956'hfffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddcddccccccccbba999888888888877788788bcddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddcdcdccaaaaaaaaabbbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd348:mariob=956'hffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddcdcccccccccbaa998888888888777887888cdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeedeeedddddddddddddddccccaaaaaaaabbaeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd349:mariob=956'hffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddcdcccccccccba998888888888877887888bcddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddccbaaaaaaabbadffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd350:mariob=956'hffffffffffffffffffffffffffffffffffffffffffddddddddddddddddddddddddcdcccccccccbbba998888888888888878889cdddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddddcdccbaaaaaaabbcffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd351:mariob=956'hffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddcdcccccccccbbba99888888888788888888bddddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddeddddddddddddddccbaaaaaabbbefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd352:mariob=956'hffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddcccccccccbbbba9988888888888888888acdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddddcdcccbaaaaabbadfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd353:mariob=956'hffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddcccccccccbcbbbba9888888888888888889cddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddddcccbaaaabcbcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd354:mariob=956'hffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddcccccccccbcbbbaa988888888888888888acddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdddddddddddddcccbaaaabbbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd355:mariob=956'hffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddcccccccccccbbbbba9988888888888888889cddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddddddddddddccccaaabbbbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd356:mariob=956'hffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddcdcccccccbbbbbbaa998888888888888889bdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddddddddcccccbaabbbbcffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd357:mariob=956'hffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddcccccccccccbbbbbbaa99888888888888888acdddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdddddddddddcdcccbaabbbbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd358:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddccccccccbbbbbbaaa98888888988888899cdddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddddcccccbabbbaefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd359:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddcccccccccccbbbbbbaaa9888888888888899bddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddcccccbabbadfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd360:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddcdcccccccccbbbbbbbbaa9988888888888899acddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddccccccbbbbbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd361:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddcdcccccccccbbbbbbbaaa9988889888888999bddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdddddddddddddcccccbbbbbeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd362:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddccccccccccbbbbbbbaaaa998888888889999acdddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeeeedededdddddddddddccccccbbbbdffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd363:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddcddccccccccccbbbbbbaaaa999888888888999acddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdddddddddddddccccccbbbbffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd364:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffeeddddddddddddddddddddddddddcccccccccbbbbbbbbaaaa99888888889999abcddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddddddcccccbbbbefffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd365:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddcccccccccbbbbbbbbaaaaa9988888888999abcddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddddccccccbbbcfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd366:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddcccccccccccbbbbbbbaaaaaa998888888999aacdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddcdccccccbbbfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd367:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddcdccccccccccbbbbbbbaaaaaa998988888999aabcdddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddddccccccbaeffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd368:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddcdcdccccccccbbbbbbaaaaaaa99988888999aabcdddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddeddddddddddddddccccccbbcffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd369:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffdddddddddddddddddddddddddddcdccccccccbbbbbbbaaaaaaa99988888999aabcddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddddddcccccccbbefffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd370:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffddddddddddddddddddddddddddddccccccccccbbbbbbbaaaaaa999988889999abbddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddddddddcccccccccbdfffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd371:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffddddddddddddddddddddddddddddcccccccccbbbbbbbaaaaaaaa99988889999abbcddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddddccccccbcfffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd372:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddcccccccccccbbbbbbaaaaaaa999a99899999abbcddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdddddddddddddcccccccbeffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd373:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddccccccccccbbbbbbaaaaaaaa99a99999999abbbddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdedddddddddddddccccccbcffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd374:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddddcccccccccbbbbbbbaaaaaaa9aa99999999abbbdddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdddddddddddddccccccbbffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd375:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddccccccccccbbbbbbaaaaaaaa99a99999999abbbddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddddddccccccaefffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd376:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddcdccccccccbbbbbbbaaaaaaa99a99999999abbbdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededdddddddddddddccccccbcfffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd377:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddddccccccccbbbbbbbbaaaaaaa99aa9999999abbbdcdddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddccccccbbeffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd378:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddccccccccccbbbbbbbbaaaaaaa9a99999999abbbdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddddcccccbdffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd379:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddcdccccccccbbbbbbbaaaaaaaa9a99999999abbbddcddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddddccccccbbffffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd380:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddcdccccccccbbbbbbbbbaaaaaa99a99999999abbbdeddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddccccccbefffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd381:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddddccccccccbbbbbbbbbaaaaaaa9aa9999999aabbcfcddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddcccccbcfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd382:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddcdccccccccbbbbbbbaaaaaaaa9aa9999999aabacfdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdededdddddddddddcccccbbfffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd383:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddddccccccccbbbbbbbbbaaaaaaa9a99999999aabacfdcddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddccccccadffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd384:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeedddddddddddddddddddddddddcdcccccccccbbbbbbbbaaaaaaa9aa9999999aabbbfecdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddddcccccbcffffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd385:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddccccccccccbbbbbbbbbaaaaaa9aa99999999abbbffcdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddddcccccbefffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd386:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffdddddddddddddddddddddddddddcccccccccccbbbbbbbaaaaaaa9aa9999999aabbbffcddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedededddddddddddddcccccbcfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd387:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddccccccccccbbbbbbbbbaaaaaa9aa99999999abbbffdcdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddccccbbfffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd388:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffddddddddddddddddddddddddddcdcccccccccbbbbbbbbbaaaaaa9aa9999999aabbbefecddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddddddddccccccbdffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd389:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffeddddddddddddddddddddddddddcccccccccccbbbbbbbabaaaaa9aa9999999aabbaeffcdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddccccbbffffffffffffffffffffffffffffffffffffffffffffffffff;
10'd390:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffedddddddddddddddddddddddddddccccccccccbbbbbbbbaaaaaa9aa99999999abbaeffdcddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddccccbefffffffffffffffffffffffffffffffffffffffffffffffff;
10'd391:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffededdddddddddddddddddddddddccccccccccbcbbbbbbbaaaaaa9aa99999999abbadffdcdddddddddddeedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddcccccadfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd392:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeddddddddddddddddddddccccccccbbbbbbbbbbaaaaaaba9999999aabbadffecdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddccccbbfffffffffffffffffffffffffffffffffffffffffffffffff;
10'd393:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeddddddddddddddccccccccccbbbbbbbbabaaaa9aa99999999aabacfffccddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddcccccbdffffffffffffffffffffffffffffffffffffffffffffffff;
10'd394:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeddddddddddddcccccccccccbbbbbbbbaaaaa9b999999999abbacfffdcdddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeeddddddddddddccccbcffffffffffffffffffffffffffffffffffffffffffffffff;
10'd395:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeedddddddddddccccccccccccbbbbbbbaaaaa9aa99999999aabbbfffeccddddddddeddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeededddddddddddccccbefffffffffffffffffffffffffffffffffffffffffffffff;
10'd396:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeedddddddddddcccccccccccbbbbbbbbbaaaa9b99a999999aabbbffffccddddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddccccbdfffffffffffffffffffffffffffffffffffffffffffffff;
10'd397:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeeeeddddddddddccccccccccbcbbbbbbabaaaaaaa9999999aabbbefffdcdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedeedddddddddddcccbbfffffffffffffffffffffffffffffffffffffffffffffff;
10'd398:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeeeeeddddddddddcccccccccccbbbbbbbbaaaaab999999999aabbbefffeccdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddccccaeffffffffffffffffffffffffffffffffffffffffffffff;
10'd399:mariob=956'hffffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeeeeeeddddddddddccccccccccccbbbbbbabaaaaaaa9999999aabbadffffccdddddddddededeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddccccbcffffffffffffffffffffffffffffffffffffffffffffff;
10'd400:mariob=956'hfffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeeeeeeedddddddddddcccccccccccbbbbbabaaaaab9a9999999aabbadffffdcdddddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddedddddddddccccbefffffffffffffffffffffffffffffffffffffffffffff;
10'd401:mariob=956'hffffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeedeeeeeedddddddddddcccccccccccbbbbbbaaaaaaaaa9a99999aabbacffffeccdddddddddddeedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddddddcccbdfffffffffffffffffffffffffffffffffffffffffffff;
10'd402:mariob=956'hfffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeeeddeeedddddddddddccccccccccccbbbbbbbbaa9abaaa999999aaabbcfffffccdddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddedddddddddcccbbfffffffffffffffffffffffffffffffffffffffffffff;
10'd403:mariob=956'hffffffffffffffffffffffffffffffffffffffeeeeeeeeeeeeeeeeeeeeeeddeedddddddddddccccccccccbcbbbbbbaaaabaaaa9a99999aabbbfffffdccdddddddddedeedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddccccbdffffffffffffffffffffffffffffffffffffffffffff;
10'd404:mariob=956'hffffffffffffffffffffffffffffffffffffffedddeeeeeeeeeeeeeeeeeeedddedddddddddccccccccccccbcbbbbbbaa9baaaaa999999aabbbeffffeccdddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddcccbcffffffffffffffffffffffffffffffffffffffffffff;
10'd405:mariob=956'hffffffffffffffffffffffffffffffeeeeffffddddddddeeeeeeeeeeeeeeeeddddddddddddddcccccccccccbbbbbbbaaabaaaaaa99999aabbbeffffeccddddddddeddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddccccbefffffffffffffffffffffffffffffffffffffffffff;
10'd406:mariob=956'hfffffffffffffffffffffffedca9888888889999abddddddeeeeeeeeeeeeeddddddddddddddccccccccccccbbbbbbbaa9bbaaaaaaa999aabbbdfffffdccdddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddddcccbcfffffffffffffffffffffffffffffffffffffffffff;
10'd407:mariob=956'hffffffffffffffffffffeca987777766676777777668acddddddeeeeeeeeedddddddddddddddccccccccccbbbbbbbbbaabaaaaaaaa999aabbbcfffffeccdddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddcccbfffffffffffffffffffffffffffffffffffffffffff;
10'd408:mariob=956'hffffffffffffffffffeb988766666666656666666666568cdddddeeeeeeeeeddddddcdddddccdccccccccbccbbbbbbaaabaaaaaaaaa99aaabbcffffffcccdddddddddeedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddcccbdffffffffffffffffffffffffffffffffffffffffff;
10'd409:mariob=956'hffffffffffffffffeb8877666665555555555555555555556addddddddeedddddddddcddddddccdcccccccbcbbbbbbbabbaaaaaaaaa99aaabbbffffffdccdddddddddedeedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddccbbffffffffffffffffffffffffffffffffffffffffff;
10'd410:mariob=956'hfffffffffffffffb98776666655555555544444444445555546acdddddddddddddddddccdddcdccccccccccbbbbbbbbabbaaaaaaaaaaaaaabbaefffffdccdddddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededddddddddddddccbefffffffffffffffffffffffffffffffffffffffff;
10'd411:mariob=956'hfffffffffffffea87766665555555544444444444444444455445addddddddddddddddddccdcccccccccccbcbbbbbbb9bbaaaaaaaaaaaaaaabadfffffecccdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddeeeeeeedddddddddbcfffffffffffffffffffffffffffffffffffffffff;
10'd412:mariob=956'hffffffffffffc977666555555544444444443333333334444444435adddddddddddddddddccdcccccccccccbcbbbbbaabaaaaaaaaaaaa99abbacffffffdccdddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddeeeeeeeeeeeeededdddddddcbeffffffffffffffffffffffffffffffffffffffff;
10'd413:mariob=956'hfffffffffffb877666555555545444444444333333333333344444336bddddddddddddddddccccccccccccccbbbbbbaabbbabaaaaaaaaaaaabbbffffffecdddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddeeeeeeeeeeeeededddddddddddbdffffffffffffffffffffffffffffffffffffffff;
10'd414:mariob=956'hffffffffffb877666555555444444444443433333333333333334444337ddcddddddddddddcccccccccccccbcbbbbbaacaabaaaaaaaaa9aaabbbefffffecdcdddddddededeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeededdddddddddddddbffffffffffffffffffffffffffffffffffffffff;
10'd415:mariob=956'hfffffffffa877666555554444444444444444333333333333333333343249ddccdddddddddddccccccccccccbcbbbbaabbbabaaaaaaaaaaaabbaeffffffdddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddddddcddcdccdcdfffffffffffffffffffffffffffffffffffffff;
10'd416:mariob=956'hffffffffb77666655555554444444444444443333333333333333333333336bccccddcddddcccccccccccccccbbbbbabbabbaaaaaaaaaa9aaabadffffffecdcdddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddddddcdcccccccccfffffffffffffffffffffffffffffffffffffff;
10'd417:mariob=956'hfffffffc87766555555544444444444444444333333333333333333333333249cccccdddcdddcccccccccccbbcbbbbabbbbabaaaaaaaaaaaaabbcffffffecddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddcddccccccbccbccccffffffffffffffffffffffffffffffffffffff;
10'd418:mariob=956'hffffffd8766665555454444445444444444444434333333333333333333333325bccccccddccddccccccccbccbbbbb9bbabbabaaaaaaaaaaaaabbfffffffdddddddddededeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddcddccccbccbbbbbbbbbcfffffffffffffffffffffffffffffffffffff;
10'd419:mariob=956'hffffff9766665555554445445555555555444444433333333333333333333333239bccccccdccccccccccccbbcbcbb9bbbbabaaaaaaaaaa9aaabbcffffffddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddddccccbccbbbabbabbaaabbbdffffffffffffffffffffffffffffffffffff;
10'd420:mariob=956'hfffffc77666555544555444555555554444454444433333332333333333333333226bcbcccccddcccccccccccbbbcbacbbababaaaaaaa9abcbbbbbefffffeddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddcccccbbbaaba9a9999899aaabbefffffffffffffffffffffffffffffffffff;
10'd421:mariob=956'hffffe87666555555544555555555555555554444433333333333233333333333333239ccccccccccccccccccccccbbaccbbbbbbbaa99accbbbbbbbbffffffddddddddedeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddccccbaaa877654554556677889aaadefffffffffffffffffffffffffffffffff;
10'd422:mariob=956'hffffb766665555554555555566666666555555444443333333322323333333333333225abcbcccccccccccccccccccabbbaaa99aabccbbbbbbbbabadfffffdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeedddddddccbba88754334445555666667778888889abdfffffffffffffffffffffffffffff;
10'd423:mariob=956'hfffe876665555554444555556666666666655554444433333332233333333333333332138bcccbccccccccccccccccbbcbbccccccbbbbbbbbbaaabacfffffdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddddcbba876433344445555555666666666777778889bdffffffffffffffffffffffffff;
10'd424:mariob=956'hfffb7666555555444555555666777776666655554443443333332233333333333333333215abbbbbcccbcccccbccccbbcccbbbbbbbbbbbaaaaaabbabfffffddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddcccba974323344444444555555555555655556666777789cffffffffffffffffffffffff;
10'd425:mariob=956'hfff9766655555454445555566777777766666655444333333333223322233333333333332137aabbbbbcbbccbcbccbcacbbbbbbbbbbbaaaa99aabbabfffffddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeddddccca98533334444444444444444444545555555556666677789cffffffffffffffffffffff;
10'd426:mariob=956'hffe776655555444454555566677777777666666555444333333332233233333333333333322149aaabbbbbbbbbbbbbbabcbbbbbbbaaaa99999aabbacfffffdddddddddeeeeeeeeeeeeeeeeeeeeeeeeeedddcccb864333444444444444444444444444444455555555565667789dffffffffffffffffffff;
10'd427:mariob=956'hffb76665555444454455556777777777877666555544443333333223232333333333333333222159aaabbabbabbbbbb9bbbbaaaaaa99999999abbbadfffffddddddddeeeeeeeeeeeeeeeeeeeeeeeeeddddcbb853234444444444444444444444444444444445555555555666778beffffffffffffffffff;
10'd428:mariob=956'hff97665555544444454555667777888777776666554433333333332222233333333333333333221269aaaaaaaaaaaaaabbaaa99999999999aaabbbbeffffedddddddeeeeeeeeeeeeeeeeeeeeeeeeddddcbb9533344444444444433433333444444444444444444555555555666779efffffffffffffffff;
10'd429:mariob=956'hfe866655555444444545665666777877777666665544433333333322323333333333333333333222136999999a9aa9a9aa9999999999999aa97abacfffffedddddddeeeeeeeeeeeeeeeeeeeeededdddcba533444444444444433433333334334444444444444444444555555666678cffffffffffffffff;
10'd430:mariob=956'hfc7665555544444445555666676778777776666654543333333333332322223333333333333333232212468999999999999999999999aa975569bbffffffdddddeddeeeeeeeeeeeeeeeeeeeddddddcba633344444444444343343333333334333444444444444444445555555566678afffffffffffffff;
10'd431:mariob=956'hfb766555554444444455566667777777777666555544433333333333322233333333333333333333333221246899999999999999998764445568acfffffeddddeeddeeeeeeeeeeeeeeeeeedddddcca843344444444444433334333333333334444444444444444444444555555556677affffffffffffff;
10'd432:mariob=956'hfa666555554444444445456566667767767666655544433333333333222223223333333333333333333333221123567788888765443334445568abfffffddddededdeeeeeeeeeeeeeeeeedddcdca963344444444444334433433333443443343444444444444444444444544555556667afffffffffffff;
10'd433:mariob=956'hf8666555544444444444555666666777666666555544433333333333322323232233333333333333333333333332222222222233333344445557aaefffeddddeeedeeeeeeeeeeeeeeeeddddccb9742344444444444433333334444443444444444444444444444444444444455555566679ffffffffffff;
10'd434:mariob=956'he8665555544444444444445566666667666655555544433333333333323333322233333333333333333333333333333333333333333434444557aadfffedddeeeedddeeeeeeeeeeeeedddccca86333444444444444333333433444444444444444444444444444444444444445555555677afffffffffff;
10'd435:mariob=956'he86655554444444444444556556666666665555444443333333333333222222333233333333333333333333333333333333333333334444445579bcfffddeddddeddeeeeeeeeeeeeedddccc97323444444444444433344444444444444444444444444444444444444444444445555556668bffffffffff;
10'd436:mariob=956'hd7665555444444444444444555555655555555544444333333333333333333322333333333333333333333333333333333333333333334444557abcffedddeeeeddeeeeeeeeeeddddddccb8422344444444444343333444444444444444544444444444444444444444444444444555556678bfffffffff;
10'd437:mariob=956'hd7665555444444444444444455555555555544444443333333333333333333333333333333333333333333333333333333333333333344444557abcffedddeeeedeeeeeeeeeedddddccba721334444444444444334433444444444444444444444444444444444444444444444444555556679cffffffff;
10'd438:mariob=956'hd7665554444444444444444444555555444454444433333333333333333333333333333333333333333333333333333333333333333334444557abcffeddeeeeedeeeeeeeeeddddcdbba4023344444444444443434444444444445455444445544444444444444444444444444444455556667adfffffff;
10'd439:mariob=956'hd7655554444444444444444444445554544444444334333333333333333333333333333333333333333333333333333333333333333334444558aacffedddeeeedeeeeeedddddcccba8202344444444444444434344444444545555555544444444444444444444444444444444444455556678aeffffff;
10'd440:mariob=956'hd7655554444444444444444444444444444444444433333333333333333333333333333333333333333333333333333333333333333334444558badfffddddeeddeeedddddddcccba501234444444444444444444444444445545555555554544444444444444444444444444444444555566679cffffff;
10'd441:mariob=956'he7655554444444443333434344444444444444443333333333333333333333333333333333333333333333333333333333333333333333444569badfffddddddeddddddddddccba82013334444444444444444444444445555555556666555544444444444444444444444444444444455556678aefffff;
10'd442:mariob=956'he865555444444443343333343444444444444343333333333333333333333333333333333333333333333333333333333333333333333444557abaefffeddddddddddddcccccb94002334444444444444444444444444555556666666666555555444444444444444444444444444444455556679bfffff;
10'd443:mariob=956'hf965555444444443333333333343444444433333333333333333333333333333333333333333333333333333333333333333333333334444558bbbfffffdcdddddddcccccbba710123344444444444444444444444555555566655666666655555544444444444444444444444444444455556668adffff;
10'd444:mariob=956'hf966555444444433333343334333444443333333333333333333333333333333333333333333333333333333333333333333333333334444569bacffffffccccccccccbcba82002333444454444444444444444444555565566667666666666555444444444444444444444444444444445555667abffff;
10'd445:mariob=956'hfb6655544444333333333333344433333333343333333333333333333333333333333333333333333333333333333333333333333344444557abbdffffffeabbccbcbbb962001233444444454444444444444444455556666666766666666655555544444444444444444444444444444445556679bdfff;
10'd446:mariob=956'hfc7655544444433333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333344445569bbbeffffffd76899a9764221223344444444554444444444444444555566666666767776776665554444444444444444444444444444444445555668acfff;
10'd447:mariob=956'hfe865554444444333333333333333333343333333333333333333333333333333333333333333333333333333333333333333333344444558bbacfffffffd8654444333333444444555455444544444444444445556566667777787777777665555444444444444443444444444444444445555667abfff;
10'd448:mariob=956'hff96655444444333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333444444557abbbefffffffd76655555554455555555555555545444444444444455556667777777778777676665554444444444444444444444444444444445556679adff;
10'd449:mariob=956'hffc665554443433333333333333333333333333333333333333333333333333333333333333333333333333333333333333333344444568abbadffffffffd76655555555555555555555555544444444444444455666667778777778777766655554444444444444444434444444444444444555678acff;
10'd450:mariob=956'hfff866555444433333333333333333333333333333333333333333333333333333333333333333333333333333333333333333444456778bbabfffffffffd86655555555555555555555555555444444444444455666667777777777776666655554444444444444444444444444444444445555568abef;
10'd451:mariob=956'hfffb76555444433333333333333333333333333333333333333333333333333333333333333333333333333333333333433334455665568bbbffffffffffe86655555555555555555555555555444444444444445566666777777777766666555444444444444444344434434444444444444555567abdf;
10'd452:mariob=956'hffff96655444433333333333333333333333333333333333333333333333333333333333333333333333333333333334444556654445568bacffffffffffe866655555555555555555555555544444444444445555666666777777776666655455444444444444443334443344444444444445555679bcf;
10'd453:mariob=956'hffffe8665544443333333333333333333333333333333333333333333333333333333333333333333333344344444555555443344455668bacfffffffffffa66655555555555555555555555544444444444444555556667676777767656555544444444444444334443343444444444444444555669bcf;
10'd454:mariob=956'hfffffe866554444333333333333333333333333333333333333333333333333333333333333333333334444455565543333444455555668bacfffffffffffb76655555555555555555555555444444444444444455555666667667666665555554444444344333333333333433444444444444555668bbf;
10'd455:mariob=956'hffffffd8665544433333333333333333333333333333333333333333333333333333333333433334444445654433334444444555555557abacfffffffffffc76655555555555555555555555444444444444444455556665566666666555554444444444434333333333333333343444444444555668bbe;
10'd456:mariob=956'hfffffffea765544444333333333333333333333333333333333333333333333333333333334344444556664334444444444555555567abbbacfffffffffffe86665555555555555555555555444444444444444445555556556655565555555444444444433433333333333333343434444444555568abe;
10'd457:mariob=956'hffffffffb8776544443333333333333333333333333333333333333333333333333333343444445565555444444444444445455679abbbbabfffffffffffffa6655555555555565555555555444444444444444445455555555555555554555444444434334333333333333333343444444444555568bbe;
10'd458:mariob=956'hffffffffb866676554433333333333333333333332333333333333333333333333333344444456554455444444444444444578abbbbbaabdffffffffffffffd7666555555555566555555555444444444444444444444555555555555454544444434344333333333333333333333444344444455668bbd;
10'd459:mariob=956'hffffffffb8776556665543333333333333333333333233333333333333333333333444445566544457754444444455678abbbbbbaaabdefffffffffffffffff9666555555655666555555554444444444444444444444455545455554444444444433333333333333333333333333344344444555568bbd;
10'd460:mariob=956'hfffffffeb887776544556554333333333333333333223333333333333333333344444555544444557bba97556789aabbbbbaaabbcdfffffffffffffffffffffb766655555666666655555554444444444444344444444444544555444444444444333333333333333333333333333333434444455568bbd;
10'd461:mariob=956'hfffffffea88877766654444455543333333333333333333333333333333333444556554444445558bbbbbbabbbbbbbaaaabcdefffffffffffffffffffffffffe976666556666666655555554444444444444433344444454444444444444444444433333333333333333333333333333334444455669bbe;
10'd462:mariob=956'hffffffffb8887777776666554444444444443333333333333333333334444555544334444555559bbbadffdbaabbbcdeffffffffffffffffffffffffffffffffc76666556666666655555544444444444433333333444444434444444444434433333333333333333333333333333333344444455679bbe;
10'd463:mariob=956'hffffffffe98777777777766666655544444444444444444444444444444444434444445555556abbbbdffffffefffffffffffffffffffffffffffffffffffffffa7665556666666655555544444444444333333333434444444444444434333333333333333333333333333333333333334444455679bbe;
10'd464:mariob=956'hffffffffffa87777777777777766666665554443333333333433333333334444444555555458bbbabeffffffffffffffffffffffffffffffffffffffffffffffff966666666666666655555444444443333333333333434444433343334434433333333333333333333333333333333334344445567abbf;
10'd465:mariob=956'hffffffffffeb98777777777777777766666666665555444444444444444444455555555568bbbbabfffffffffffffffffffffffffffffffffffffffffffffffffff97666666666666655554444444444433333333333333333444334434333333333333333333333333333333333333333444445568abbf;
10'd466:mariob=956'hffffffffffffcba987777777777777777666666666666555555444444455555555555569abbbabdffffffffffffffffffffffffffffffffffffffffffffffffffffa8776666666666665555444444444333333333333333333343444433333333333333333333333333333333333333333444455568bacf;
10'd467:mariob=956'hffffffffffffffdbaaa98766777777777666666666666666666555555555555444568abbbbaacffffffffffffffffffffffffffffffffffffffffffffffffffffffb7677766666676665555444444433333333333333333343333333333333333333333333333333333333333333333334444455579bacf;
10'd468:mariob=956'hfffffffffffffffffdbbbba9877666666766666666666666666665555554445679bbbbbaabdffffffffffffffffffffffffffffffffffffffffffffffffffffffffb8755787767777665555544444444333333333333333333333333333333333333333333333333333333333333333333444455679badf;
10'd469:mariob=956'hffffffffffffffffffffdcbbbaaa9877666666666666666655555555556789abbbbbaabceffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb887655787777766655554444433433333333333333333333333333333333333333333333333333333333333333333344445568abbef;
10'd470:mariob=956'hfffffffffffffffffffffffedcbaabbbbaaa99988777777667778899aabbbbbbaaabdefffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc887765457877766655554444444333333333333333333333333333333333333333333333333333333333333333333444455668bbbff;
10'd471:mariob=956'hffffffffffffffffffffffffffffedccbbbaabbbbbbbbbbbbbbbbbbbbbaaabbcdeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb8777765457877665555444443443333333333333333333333333333333333333333333333333333333333333333334445566abacff;
10'd472:mariob=956'hfffffffffffffffffffffffffffffffffffeddcccbbbbbbbbbbbbbbbccddeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb877776555688766555544444343333333333333333333333333333333333333333333333333333333333333333334445567bbadff;
10'd473:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc87777655458876555544444443333333333333333333333333333333333333333333333333333333333333333444455679bbbfff;
10'd474:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda97777653498665555444434333333333333333333333333333333333333333333333333333333333333333344445568abacfff;
10'd475:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeca98776338a765555444443433333333333333333333333333333333333333333333333333333333333333344455579bbbdfff;
10'd476:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecba98436a97655554444433333333333333333333333333333333333333333333333333333333333333344445568bbacffff;
10'd477:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcbbaaba8886654444444333333333333333333333333333333333333333333333333333333333333444445567abbbeffff;
10'd478:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbaa9888655544444333333333333333333333333333333333333333333333333333333333334444445579bbacfffff;
10'd479:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffec997786554444443333333333333333333333333333333333333333333333333333333333344445569bbabffffff;
10'd480:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb9877776554444433333333333333333333333333333333333333333333333333333333444455669bbbbeffffff;
10'd481:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd988767765444443333333333333333333333333333333333333333333333333333344344455679bbbadfffffff;
10'd482:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc888766776544433333333333333333333333333332333333333333333333333334444445669abbbadffffffff;
10'd483:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa8877655666544333333333333333333333333333333333333333333333333444444556778bbbabdfffffffff;
10'd484:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe9887766556665444333333333333333333333333333333333333333333344444455676668bbabeffffffffff;
10'd485:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd877777665455655443333333333333233333332333333333333333444444556666555678bbaefffffffffff;
10'd486:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd87777766654445555443333333333333333333333333333334444455566655444555678bbaefffffffffff;
10'd487:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd8777777666654444455554443333333333333333333444455566665544334455556678bbaefffffffffff;
10'd488:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd877777766666655443334455555554444455555556555554433333444445555566679bbaefffffffffff;
10'd489:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffea777777776666666555443333334444444443333333333334444444555555556668abbbffffffffffff;
10'd490:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffb8767777766666666666555544433333344444444444444444555555555555667abbacffffffffffff;
10'd491:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffda8766777676666666666666666555544444444444555555555555555555579bbbabfffffffffffff;
10'd492:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffcb977666766777666666666666666666555555555555555555555555679bbbbabffffffffffffff;
10'd493:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecba976666666676666666666666666666666555555555555555679abbbaabdfffffffffffffff;
10'd494:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdbbba8776666666666666666666666666666665554556789bbbbbaaabdfffffffffffffffff;
10'd495:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffecbbaaa987666666666666666665665666667789aabbbbbaaabcdffffffffffffffffffff;
10'd496:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffedcbabbbaa9988776666677888999aaabbbbbbbaaaabcdefffffffffffffffffffffff;
10'd497:mariob=956'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffdccbbabbbbbbbbbbbbbbbbbbbbaaaaabbccdeffffffffffffffffffffffffffff;
10'd498:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeddcbbbbbbbbbbbbbbcccddeefffffffffffffffffffffffffffffffffff;
10'd499:mariob=956'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;


	endcase
end				
						
						
endmodule











