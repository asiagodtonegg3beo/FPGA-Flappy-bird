module state(ix_index,iy_index,imode,clk);
input ix_index;
input iy_index;
input imode;
input clk;

parameter air = 4'h0,question = 4'h1,coin = 4'h2;
parameter w_length = 844;
reg [w_length-1:0] map;

always@(posedge clk)
begin

case(iy_index)
4'h0:map = 844'h000000000000000000000000000000000000000000000000000;
4'h1:map = 844'h000000000000000000000000000000000000000000000000000;
4'h2:map = 844'h000000000000002000000000000000000000000000000000000;
4'h3:map = 844'h000000000000001000000000000000000000000000000000000;
4'h4:map = 844'h000000000000000000000000000000000000000000000000000;
4'h5:map = 844'h000000000000000000000000000000000000000000000000000;
4'h6:map = 844'h000000000000022200000000000000000000000000000000000;
4'h7:map = 844'h000000001000010100000000000000000000000000000000000;
4'h8:map = 844'h000000000000000000000000000000000000000000000000000;
4'h9:map = 844'h000000000000000000000000000000000000000000000000000;
4'ha:map = 844'h000000000000000000000000000000000000000000000000000;
4'hb:map = 844'h000000000000000000000000000000000000000000000000000;
4'hc:map = 844'h000000000000000000000000000000000000000000000000000;
endcase

end

endmodule